-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity initialiseCounters is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(1 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity initialiseCounters;
architecture initialiseCounters_arch of initialiseCounters is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal initialiseCounters_CP_3_start: Boolean;
  signal initialiseCounters_CP_3_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal if_stmt_98_branch_ack_1 : boolean;
  signal if_stmt_98_branch_ack_0 : boolean;
  signal array_obj_ref_95_index_0_scale_req_0 : boolean;
  signal array_obj_ref_95_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_95_index_0_scale_req_1 : boolean;
  signal array_obj_ref_95_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_95_index_sum_1_req_0 : boolean;
  signal array_obj_ref_95_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_95_index_sum_1_req_1 : boolean;
  signal array_obj_ref_95_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_95_store_0_req_0 : boolean;
  signal array_obj_ref_95_store_0_ack_0 : boolean;
  signal array_obj_ref_95_store_0_req_1 : boolean;
  signal array_obj_ref_95_store_0_ack_1 : boolean;
  signal if_stmt_98_branch_req_0 : boolean;
  signal phi_stmt_82_req_0 : boolean;
  signal nJ_92_86_buf_req_0 : boolean;
  signal nJ_92_86_buf_ack_0 : boolean;
  signal nJ_92_86_buf_req_1 : boolean;
  signal nJ_92_86_buf_ack_1 : boolean;
  signal phi_stmt_82_req_1 : boolean;
  signal phi_stmt_82_ack_0 : boolean;
  signal if_stmt_105_branch_req_0 : boolean;
  signal if_stmt_105_branch_ack_1 : boolean;
  signal if_stmt_105_branch_ack_0 : boolean;
  signal phi_stmt_69_req_0 : boolean;
  signal nI_79_73_buf_req_0 : boolean;
  signal nI_79_73_buf_ack_0 : boolean;
  signal nI_79_73_buf_req_1 : boolean;
  signal nI_79_73_buf_ack_1 : boolean;
  signal phi_stmt_69_req_1 : boolean;
  signal phi_stmt_69_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "initialiseCounters_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  initialiseCounters_CP_3_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "initialiseCounters_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= initialiseCounters_CP_3_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= initialiseCounters_CP_3_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= initialiseCounters_CP_3_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  initialiseCounters_CP_3: Block -- control-path 
    signal initialiseCounters_CP_3_elements: BooleanArray(24 downto 0);
    -- 
  begin -- 
    initialiseCounters_CP_3_elements(0) <= initialiseCounters_CP_3_start;
    initialiseCounters_CP_3_symbol <= initialiseCounters_CP_3_elements(18);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	19 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_67/$entry
      -- CP-element group 0: 	 branch_block_stmt_67/branch_block_stmt_67__entry__
      -- CP-element group 0: 	 branch_block_stmt_67/merge_stmt_68__entry__
      -- CP-element group 0: 	 branch_block_stmt_67/merge_stmt_68_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_67/merge_stmt_68__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_67/merge_stmt_68__entry___PhiReq/phi_stmt_69/$entry
      -- CP-element group 0: 	 branch_block_stmt_67/merge_stmt_68__entry___PhiReq/phi_stmt_69/phi_stmt_69_sources/$entry
      -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	16 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	8 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_scale_0_sample_complete
      -- CP-element group 1: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_scale_0_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_scale_0_Sample/ra
      -- 
    ra_59_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_95_index_0_scale_ack_0, ack => initialiseCounters_CP_3_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	16 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (4) 
      -- CP-element group 2: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_scaled_0
      -- CP-element group 2: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_scale_0_update_complete
      -- CP-element group 2: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_scale_0_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_scale_0_Update/ca
      -- 
    ca_64_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_95_index_0_scale_ack_1, ack => initialiseCounters_CP_3_elements(2)); -- 
    -- CP-element group 3:  join  transition  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: 	16 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_partial_sum_1_sample_start
      -- CP-element group 3: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_partial_sum_1_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_partial_sum_1_Sample/rr
      -- 
    rr_85_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_85_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialiseCounters_CP_3_elements(3), ack => array_obj_ref_95_index_sum_1_req_0); -- 
    initialiseCounters_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "initialiseCounters_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initialiseCounters_CP_3_elements(2) & initialiseCounters_CP_3_elements(16);
      gj_initialiseCounters_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initialiseCounters_CP_3_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	8 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_partial_sum_1_sample_complete
      -- CP-element group 4: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_partial_sum_1_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_partial_sum_1_Sample/ra
      -- 
    ra_86_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_95_index_sum_1_ack_0, ack => initialiseCounters_CP_3_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	16 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (27) 
      -- CP-element group 5: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_offset_calculated
      -- CP-element group 5: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_word_address_calculated
      -- CP-element group 5: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_root_address_calculated
      -- CP-element group 5: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_partial_sum_1_update_complete
      -- CP-element group 5: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_partial_sum_1_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_partial_sum_1_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_final_index_sum_regn/$entry
      -- CP-element group 5: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_final_index_sum_regn/$exit
      -- CP-element group 5: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_final_index_sum_regn/req
      -- CP-element group 5: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_final_index_sum_regn/ack
      -- CP-element group 5: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_base_plus_offset/$entry
      -- CP-element group 5: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_base_plus_offset/$exit
      -- CP-element group 5: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_base_plus_offset/sum_rename_req
      -- CP-element group 5: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_base_plus_offset/sum_rename_ack
      -- CP-element group 5: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_word_addrgen/$entry
      -- CP-element group 5: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_word_addrgen/$exit
      -- CP-element group 5: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_word_addrgen/root_register_req
      -- CP-element group 5: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_word_addrgen/root_register_ack
      -- CP-element group 5: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_Sample/array_obj_ref_95_Split/$entry
      -- CP-element group 5: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_Sample/array_obj_ref_95_Split/$exit
      -- CP-element group 5: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_Sample/array_obj_ref_95_Split/split_req
      -- CP-element group 5: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_Sample/array_obj_ref_95_Split/split_ack
      -- CP-element group 5: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_Sample/word_access_start/$entry
      -- CP-element group 5: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_Sample/word_access_start/word_0/$entry
      -- CP-element group 5: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_Sample/word_access_start/word_0/rr
      -- 
    ca_91_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_95_index_sum_1_ack_1, ack => initialiseCounters_CP_3_elements(5)); -- 
    rr_121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialiseCounters_CP_3_elements(5), ack => array_obj_ref_95_store_0_req_0); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (5) 
      -- CP-element group 6: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_Sample/word_access_start/$exit
      -- CP-element group 6: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_Sample/word_access_start/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_Sample/word_access_start/word_0/ra
      -- 
    ra_122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_95_store_0_ack_0, ack => initialiseCounters_CP_3_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	16 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_Update/word_access_complete/$exit
      -- CP-element group 7: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_Update/word_access_complete/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_Update/word_access_complete/word_0/ca
      -- 
    ca_133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_95_store_0_ack_1, ack => initialiseCounters_CP_3_elements(7)); -- 
    -- CP-element group 8:  branch  join  transition  place  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	1 
    -- CP-element group 8: 	4 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	10 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (24) 
      -- CP-element group 8: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97__exit__
      -- CP-element group 8: 	 branch_block_stmt_67/branch_block_stmt_80/if_stmt_98__entry__
      -- CP-element group 8: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/$exit
      -- CP-element group 8: 	 branch_block_stmt_67/branch_block_stmt_80/ULT_u8_u1_101_place
      -- CP-element group 8: 	 branch_block_stmt_67/branch_block_stmt_80/if_stmt_98_if_link/$entry
      -- CP-element group 8: 	 branch_block_stmt_67/branch_block_stmt_80/if_stmt_98_else_link/$entry
      -- CP-element group 8: 	 branch_block_stmt_67/branch_block_stmt_80/if_stmt_98_dead_link/$entry
      -- CP-element group 8: 	 branch_block_stmt_67/branch_block_stmt_80/if_stmt_98_eval_test/$entry
      -- CP-element group 8: 	 branch_block_stmt_67/branch_block_stmt_80/if_stmt_98_eval_test/$exit
      -- CP-element group 8: 	 branch_block_stmt_67/branch_block_stmt_80/if_stmt_98_eval_test/ULT_u8_u1_101/$entry
      -- CP-element group 8: 	 branch_block_stmt_67/branch_block_stmt_80/if_stmt_98_eval_test/ULT_u8_u1_101/$exit
      -- CP-element group 8: 	 branch_block_stmt_67/branch_block_stmt_80/if_stmt_98_eval_test/ULT_u8_u1_101/ULT_u8_u1_101_inputs/$entry
      -- CP-element group 8: 	 branch_block_stmt_67/branch_block_stmt_80/if_stmt_98_eval_test/ULT_u8_u1_101/ULT_u8_u1_101_inputs/$exit
      -- CP-element group 8: 	 branch_block_stmt_67/branch_block_stmt_80/if_stmt_98_eval_test/ULT_u8_u1_101/SplitProtocol/$entry
      -- CP-element group 8: 	 branch_block_stmt_67/branch_block_stmt_80/if_stmt_98_eval_test/ULT_u8_u1_101/SplitProtocol/$exit
      -- CP-element group 8: 	 branch_block_stmt_67/branch_block_stmt_80/if_stmt_98_eval_test/ULT_u8_u1_101/SplitProtocol/Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_67/branch_block_stmt_80/if_stmt_98_eval_test/ULT_u8_u1_101/SplitProtocol/Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_67/branch_block_stmt_80/if_stmt_98_eval_test/ULT_u8_u1_101/SplitProtocol/Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_67/branch_block_stmt_80/if_stmt_98_eval_test/ULT_u8_u1_101/SplitProtocol/Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_67/branch_block_stmt_80/if_stmt_98_eval_test/ULT_u8_u1_101/SplitProtocol/Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_67/branch_block_stmt_80/if_stmt_98_eval_test/ULT_u8_u1_101/SplitProtocol/Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_67/branch_block_stmt_80/if_stmt_98_eval_test/ULT_u8_u1_101/SplitProtocol/Update/cr
      -- CP-element group 8: 	 branch_block_stmt_67/branch_block_stmt_80/if_stmt_98_eval_test/ULT_u8_u1_101/SplitProtocol/Update/ca
      -- CP-element group 8: 	 branch_block_stmt_67/branch_block_stmt_80/if_stmt_98_eval_test/branch_req
      -- 
    branch_req_160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialiseCounters_CP_3_elements(8), ack => if_stmt_98_branch_req_0); -- 
    initialiseCounters_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "initialiseCounters_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initialiseCounters_CP_3_elements(1) & initialiseCounters_CP_3_elements(4) & initialiseCounters_CP_3_elements(7);
      gj_initialiseCounters_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initialiseCounters_CP_3_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  fork  transition  place  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	13 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (11) 
      -- CP-element group 9: 	 branch_block_stmt_67/branch_block_stmt_80/if_stmt_98_if_link/$exit
      -- CP-element group 9: 	 branch_block_stmt_67/branch_block_stmt_80/if_stmt_98_if_link/if_choice_transition
      -- CP-element group 9: 	 branch_block_stmt_67/branch_block_stmt_80/J_loopback
      -- CP-element group 9: 	 branch_block_stmt_67/branch_block_stmt_80/J_loopback_PhiReq/$entry
      -- CP-element group 9: 	 branch_block_stmt_67/branch_block_stmt_80/J_loopback_PhiReq/phi_stmt_82/$entry
      -- CP-element group 9: 	 branch_block_stmt_67/branch_block_stmt_80/J_loopback_PhiReq/phi_stmt_82/phi_stmt_82_sources/$entry
      -- CP-element group 9: 	 branch_block_stmt_67/branch_block_stmt_80/J_loopback_PhiReq/phi_stmt_82/phi_stmt_82_sources/Interlock/$entry
      -- CP-element group 9: 	 branch_block_stmt_67/branch_block_stmt_80/J_loopback_PhiReq/phi_stmt_82/phi_stmt_82_sources/Interlock/Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_67/branch_block_stmt_80/J_loopback_PhiReq/phi_stmt_82/phi_stmt_82_sources/Interlock/Sample/req
      -- CP-element group 9: 	 branch_block_stmt_67/branch_block_stmt_80/J_loopback_PhiReq/phi_stmt_82/phi_stmt_82_sources/Interlock/Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_67/branch_block_stmt_80/J_loopback_PhiReq/phi_stmt_82/phi_stmt_82_sources/Interlock/Update/req
      -- 
    if_choice_transition_165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_98_branch_ack_1, ack => initialiseCounters_CP_3_elements(9)); -- 
    req_201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialiseCounters_CP_3_elements(9), ack => nJ_92_86_buf_req_0); -- 
    req_206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialiseCounters_CP_3_elements(9), ack => nJ_92_86_buf_req_1); -- 
    -- CP-element group 10:  merge  branch  transition  place  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	8 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	18 
    -- CP-element group 10: 	17 
    -- CP-element group 10:  members (28) 
      -- CP-element group 10: 	 branch_block_stmt_67/branch_block_stmt_80__exit__
      -- CP-element group 10: 	 branch_block_stmt_67/if_stmt_105__entry__
      -- CP-element group 10: 	 branch_block_stmt_67/branch_block_stmt_80/$exit
      -- CP-element group 10: 	 branch_block_stmt_67/branch_block_stmt_80/branch_block_stmt_80__exit__
      -- CP-element group 10: 	 branch_block_stmt_67/branch_block_stmt_80/if_stmt_98__exit__
      -- CP-element group 10: 	 branch_block_stmt_67/branch_block_stmt_80/if_stmt_98_else_link/$exit
      -- CP-element group 10: 	 branch_block_stmt_67/branch_block_stmt_80/if_stmt_98_else_link/else_choice_transition
      -- CP-element group 10: 	 branch_block_stmt_67/if_stmt_105_dead_link/$entry
      -- CP-element group 10: 	 branch_block_stmt_67/if_stmt_105_eval_test/$entry
      -- CP-element group 10: 	 branch_block_stmt_67/if_stmt_105_eval_test/$exit
      -- CP-element group 10: 	 branch_block_stmt_67/if_stmt_105_eval_test/ULT_u8_u1_108/$entry
      -- CP-element group 10: 	 branch_block_stmt_67/if_stmt_105_eval_test/ULT_u8_u1_108/$exit
      -- CP-element group 10: 	 branch_block_stmt_67/if_stmt_105_eval_test/ULT_u8_u1_108/ULT_u8_u1_108_inputs/$entry
      -- CP-element group 10: 	 branch_block_stmt_67/if_stmt_105_eval_test/ULT_u8_u1_108/ULT_u8_u1_108_inputs/$exit
      -- CP-element group 10: 	 branch_block_stmt_67/if_stmt_105_eval_test/ULT_u8_u1_108/SplitProtocol/$entry
      -- CP-element group 10: 	 branch_block_stmt_67/if_stmt_105_eval_test/ULT_u8_u1_108/SplitProtocol/$exit
      -- CP-element group 10: 	 branch_block_stmt_67/if_stmt_105_eval_test/ULT_u8_u1_108/SplitProtocol/Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_67/if_stmt_105_eval_test/ULT_u8_u1_108/SplitProtocol/Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_67/if_stmt_105_eval_test/ULT_u8_u1_108/SplitProtocol/Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_67/if_stmt_105_eval_test/ULT_u8_u1_108/SplitProtocol/Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_67/if_stmt_105_eval_test/ULT_u8_u1_108/SplitProtocol/Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_67/if_stmt_105_eval_test/ULT_u8_u1_108/SplitProtocol/Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_67/if_stmt_105_eval_test/ULT_u8_u1_108/SplitProtocol/Update/cr
      -- CP-element group 10: 	 branch_block_stmt_67/if_stmt_105_eval_test/ULT_u8_u1_108/SplitProtocol/Update/ca
      -- CP-element group 10: 	 branch_block_stmt_67/if_stmt_105_eval_test/branch_req
      -- CP-element group 10: 	 branch_block_stmt_67/ULT_u8_u1_108_place
      -- CP-element group 10: 	 branch_block_stmt_67/if_stmt_105_if_link/$entry
      -- CP-element group 10: 	 branch_block_stmt_67/if_stmt_105_else_link/$entry
      -- 
    else_choice_transition_169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_98_branch_ack_0, ack => initialiseCounters_CP_3_elements(10)); -- 
    branch_req_240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialiseCounters_CP_3_elements(10), ack => if_stmt_105_branch_req_0); -- 
    -- CP-element group 11:  transition  output  delay-element  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	24 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	15 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_67/branch_block_stmt_80/merge_stmt_81__entry___PhiReq/$exit
      -- CP-element group 11: 	 branch_block_stmt_67/branch_block_stmt_80/merge_stmt_81__entry___PhiReq/phi_stmt_82/$exit
      -- CP-element group 11: 	 branch_block_stmt_67/branch_block_stmt_80/merge_stmt_81__entry___PhiReq/phi_stmt_82/phi_stmt_82_sources/$exit
      -- CP-element group 11: 	 branch_block_stmt_67/branch_block_stmt_80/merge_stmt_81__entry___PhiReq/phi_stmt_82/phi_stmt_82_sources/type_cast_85_konst_delay_trans
      -- CP-element group 11: 	 branch_block_stmt_67/branch_block_stmt_80/merge_stmt_81__entry___PhiReq/phi_stmt_82/phi_stmt_82_req
      -- 
    phi_stmt_82_req_185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_82_req_185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialiseCounters_CP_3_elements(11), ack => phi_stmt_82_req_0); -- 
    -- Element group initialiseCounters_CP_3_elements(11) is a control-delay.
    cp_element_11_delay: control_delay_element  generic map(name => " 11_delay", delay_value => 1)  port map(req => initialiseCounters_CP_3_elements(24), ack => initialiseCounters_CP_3_elements(11), clk => clk, reset =>reset);
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (2) 
      -- CP-element group 12: 	 branch_block_stmt_67/branch_block_stmt_80/J_loopback_PhiReq/phi_stmt_82/phi_stmt_82_sources/Interlock/Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_67/branch_block_stmt_80/J_loopback_PhiReq/phi_stmt_82/phi_stmt_82_sources/Interlock/Sample/ack
      -- 
    ack_202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nJ_92_86_buf_ack_0, ack => initialiseCounters_CP_3_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_67/branch_block_stmt_80/J_loopback_PhiReq/phi_stmt_82/phi_stmt_82_sources/Interlock/Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_67/branch_block_stmt_80/J_loopback_PhiReq/phi_stmt_82/phi_stmt_82_sources/Interlock/Update/ack
      -- 
    ack_207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nJ_92_86_buf_ack_1, ack => initialiseCounters_CP_3_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (5) 
      -- CP-element group 14: 	 branch_block_stmt_67/branch_block_stmt_80/J_loopback_PhiReq/$exit
      -- CP-element group 14: 	 branch_block_stmt_67/branch_block_stmt_80/J_loopback_PhiReq/phi_stmt_82/$exit
      -- CP-element group 14: 	 branch_block_stmt_67/branch_block_stmt_80/J_loopback_PhiReq/phi_stmt_82/phi_stmt_82_sources/$exit
      -- CP-element group 14: 	 branch_block_stmt_67/branch_block_stmt_80/J_loopback_PhiReq/phi_stmt_82/phi_stmt_82_sources/Interlock/$exit
      -- CP-element group 14: 	 branch_block_stmt_67/branch_block_stmt_80/J_loopback_PhiReq/phi_stmt_82/phi_stmt_82_req
      -- 
    phi_stmt_82_req_208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_82_req_208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialiseCounters_CP_3_elements(14), ack => phi_stmt_82_req_1); -- 
    initialiseCounters_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "initialiseCounters_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initialiseCounters_CP_3_elements(13) & initialiseCounters_CP_3_elements(12);
      gj_initialiseCounters_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initialiseCounters_CP_3_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  merge  transition  place  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	11 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (2) 
      -- CP-element group 15: 	 branch_block_stmt_67/branch_block_stmt_80/merge_stmt_81_PhiReqMerge
      -- CP-element group 15: 	 branch_block_stmt_67/branch_block_stmt_80/merge_stmt_81_PhiAck/$entry
      -- 
    initialiseCounters_CP_3_elements(15) <= OrReduce(initialiseCounters_CP_3_elements(11) & initialiseCounters_CP_3_elements(14));
    -- CP-element group 16:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: 	3 
    -- CP-element group 16: 	1 
    -- CP-element group 16: 	7 
    -- CP-element group 16: 	5 
    -- CP-element group 16:  members (36) 
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_resized_0
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_computed_0
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/merge_stmt_81__exit__
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97__entry__
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/$entry
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_update_start_
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_resize_0/$entry
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_resize_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_resize_0/index_resize_req
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_resize_0/index_resize_ack
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_scale_0_sample_start
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_scale_0_update_start
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_scale_0_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_scale_0_Sample/rr
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_scale_0_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_scale_0_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_resized_1
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_scaled_1
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_computed_1
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_resize_1/$entry
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_resize_1/$exit
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_resize_1/index_resize_req
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_resize_1/index_resize_ack
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_scale_1/$entry
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_scale_1/$exit
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_scale_1/scale_rename_req
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_index_scale_1/scale_rename_ack
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_partial_sum_1_update_start
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_partial_sum_1_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_partial_sum_1_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_Update/word_access_complete/$entry
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_Update/word_access_complete/word_0/$entry
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/assign_stmt_92_to_assign_stmt_97/array_obj_ref_95_Update/word_access_complete/word_0/cr
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/merge_stmt_81_PhiAck/$exit
      -- CP-element group 16: 	 branch_block_stmt_67/branch_block_stmt_80/merge_stmt_81_PhiAck/phi_stmt_82_ack
      -- 
    phi_stmt_82_ack_213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_82_ack_0, ack => initialiseCounters_CP_3_elements(16)); -- 
    rr_58_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_58_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialiseCounters_CP_3_elements(16), ack => array_obj_ref_95_index_0_scale_req_0); -- 
    cr_63_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_63_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialiseCounters_CP_3_elements(16), ack => array_obj_ref_95_index_0_scale_req_1); -- 
    cr_90_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_90_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialiseCounters_CP_3_elements(16), ack => array_obj_ref_95_index_sum_1_req_1); -- 
    cr_132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialiseCounters_CP_3_elements(16), ack => array_obj_ref_95_store_0_req_1); -- 
    -- CP-element group 17:  fork  transition  place  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	10 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	20 
    -- CP-element group 17: 	21 
    -- CP-element group 17:  members (11) 
      -- CP-element group 17: 	 branch_block_stmt_67/if_stmt_105_if_link/$exit
      -- CP-element group 17: 	 branch_block_stmt_67/if_stmt_105_if_link/if_choice_transition
      -- CP-element group 17: 	 branch_block_stmt_67/I_loopback
      -- CP-element group 17: 	 branch_block_stmt_67/I_loopback_PhiReq/$entry
      -- CP-element group 17: 	 branch_block_stmt_67/I_loopback_PhiReq/phi_stmt_69/$entry
      -- CP-element group 17: 	 branch_block_stmt_67/I_loopback_PhiReq/phi_stmt_69/phi_stmt_69_sources/$entry
      -- CP-element group 17: 	 branch_block_stmt_67/I_loopback_PhiReq/phi_stmt_69/phi_stmt_69_sources/Interlock/$entry
      -- CP-element group 17: 	 branch_block_stmt_67/I_loopback_PhiReq/phi_stmt_69/phi_stmt_69_sources/Interlock/Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_67/I_loopback_PhiReq/phi_stmt_69/phi_stmt_69_sources/Interlock/Sample/req
      -- CP-element group 17: 	 branch_block_stmt_67/I_loopback_PhiReq/phi_stmt_69/phi_stmt_69_sources/Interlock/Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_67/I_loopback_PhiReq/phi_stmt_69/phi_stmt_69_sources/Interlock/Update/req
      -- 
    if_choice_transition_245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_105_branch_ack_1, ack => initialiseCounters_CP_3_elements(17)); -- 
    req_281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialiseCounters_CP_3_elements(17), ack => nI_79_73_buf_req_0); -- 
    req_286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialiseCounters_CP_3_elements(17), ack => nI_79_73_buf_req_1); -- 
    -- CP-element group 18:  merge  transition  place  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	10 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 $exit
      -- CP-element group 18: 	 branch_block_stmt_67/$exit
      -- CP-element group 18: 	 branch_block_stmt_67/branch_block_stmt_67__exit__
      -- CP-element group 18: 	 branch_block_stmt_67/if_stmt_105__exit__
      -- CP-element group 18: 	 branch_block_stmt_67/if_stmt_105_else_link/$exit
      -- CP-element group 18: 	 branch_block_stmt_67/if_stmt_105_else_link/else_choice_transition
      -- 
    else_choice_transition_249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_105_branch_ack_0, ack => initialiseCounters_CP_3_elements(18)); -- 
    -- CP-element group 19:  transition  output  delay-element  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	0 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	23 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_67/merge_stmt_68__entry___PhiReq/$exit
      -- CP-element group 19: 	 branch_block_stmt_67/merge_stmt_68__entry___PhiReq/phi_stmt_69/$exit
      -- CP-element group 19: 	 branch_block_stmt_67/merge_stmt_68__entry___PhiReq/phi_stmt_69/phi_stmt_69_sources/$exit
      -- CP-element group 19: 	 branch_block_stmt_67/merge_stmt_68__entry___PhiReq/phi_stmt_69/phi_stmt_69_sources/type_cast_72_konst_delay_trans
      -- CP-element group 19: 	 branch_block_stmt_67/merge_stmt_68__entry___PhiReq/phi_stmt_69/phi_stmt_69_req
      -- 
    phi_stmt_69_req_265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_69_req_265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialiseCounters_CP_3_elements(19), ack => phi_stmt_69_req_0); -- 
    -- Element group initialiseCounters_CP_3_elements(19) is a control-delay.
    cp_element_19_delay: control_delay_element  generic map(name => " 19_delay", delay_value => 1)  port map(req => initialiseCounters_CP_3_elements(0), ack => initialiseCounters_CP_3_elements(19), clk => clk, reset =>reset);
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	17 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	22 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_67/I_loopback_PhiReq/phi_stmt_69/phi_stmt_69_sources/Interlock/Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_67/I_loopback_PhiReq/phi_stmt_69/phi_stmt_69_sources/Interlock/Sample/ack
      -- 
    ack_282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nI_79_73_buf_ack_0, ack => initialiseCounters_CP_3_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	17 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_67/I_loopback_PhiReq/phi_stmt_69/phi_stmt_69_sources/Interlock/Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_67/I_loopback_PhiReq/phi_stmt_69/phi_stmt_69_sources/Interlock/Update/ack
      -- 
    ack_287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nI_79_73_buf_ack_1, ack => initialiseCounters_CP_3_elements(21)); -- 
    -- CP-element group 22:  join  transition  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (5) 
      -- CP-element group 22: 	 branch_block_stmt_67/I_loopback_PhiReq/$exit
      -- CP-element group 22: 	 branch_block_stmt_67/I_loopback_PhiReq/phi_stmt_69/$exit
      -- CP-element group 22: 	 branch_block_stmt_67/I_loopback_PhiReq/phi_stmt_69/phi_stmt_69_sources/$exit
      -- CP-element group 22: 	 branch_block_stmt_67/I_loopback_PhiReq/phi_stmt_69/phi_stmt_69_sources/Interlock/$exit
      -- CP-element group 22: 	 branch_block_stmt_67/I_loopback_PhiReq/phi_stmt_69/phi_stmt_69_req
      -- 
    phi_stmt_69_req_288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_69_req_288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialiseCounters_CP_3_elements(22), ack => phi_stmt_69_req_1); -- 
    initialiseCounters_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "initialiseCounters_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initialiseCounters_CP_3_elements(20) & initialiseCounters_CP_3_elements(21);
      gj_initialiseCounters_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initialiseCounters_CP_3_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  merge  transition  place  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	19 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_67/merge_stmt_68_PhiReqMerge
      -- CP-element group 23: 	 branch_block_stmt_67/merge_stmt_68_PhiAck/$entry
      -- 
    initialiseCounters_CP_3_elements(23) <= OrReduce(initialiseCounters_CP_3_elements(19) & initialiseCounters_CP_3_elements(22));
    -- CP-element group 24:  merge  branch  transition  place  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	11 
    -- CP-element group 24:  members (15) 
      -- CP-element group 24: 	 branch_block_stmt_67/merge_stmt_68__exit__
      -- CP-element group 24: 	 branch_block_stmt_67/assign_stmt_79__entry__
      -- CP-element group 24: 	 branch_block_stmt_67/assign_stmt_79__exit__
      -- CP-element group 24: 	 branch_block_stmt_67/branch_block_stmt_80__entry__
      -- CP-element group 24: 	 branch_block_stmt_67/assign_stmt_79/$entry
      -- CP-element group 24: 	 branch_block_stmt_67/assign_stmt_79/$exit
      -- CP-element group 24: 	 branch_block_stmt_67/branch_block_stmt_80/$entry
      -- CP-element group 24: 	 branch_block_stmt_67/branch_block_stmt_80/branch_block_stmt_80__entry__
      -- CP-element group 24: 	 branch_block_stmt_67/branch_block_stmt_80/merge_stmt_81__entry__
      -- CP-element group 24: 	 branch_block_stmt_67/branch_block_stmt_80/merge_stmt_81_dead_link/$entry
      -- CP-element group 24: 	 branch_block_stmt_67/branch_block_stmt_80/merge_stmt_81__entry___PhiReq/$entry
      -- CP-element group 24: 	 branch_block_stmt_67/branch_block_stmt_80/merge_stmt_81__entry___PhiReq/phi_stmt_82/$entry
      -- CP-element group 24: 	 branch_block_stmt_67/branch_block_stmt_80/merge_stmt_81__entry___PhiReq/phi_stmt_82/phi_stmt_82_sources/$entry
      -- CP-element group 24: 	 branch_block_stmt_67/merge_stmt_68_PhiAck/$exit
      -- CP-element group 24: 	 branch_block_stmt_67/merge_stmt_68_PhiAck/phi_stmt_69_ack
      -- 
    phi_stmt_69_ack_293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_69_ack_0, ack => initialiseCounters_CP_3_elements(24)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal I_69 : std_logic_vector(7 downto 0);
    signal J_82 : std_logic_vector(7 downto 0);
    signal R_I_93_resized : std_logic_vector(3 downto 0);
    signal R_I_93_scaled : std_logic_vector(3 downto 0);
    signal R_J_94_resized : std_logic_vector(3 downto 0);
    signal R_J_94_scaled : std_logic_vector(3 downto 0);
    signal R_ZERO_2_96_wire_constant : std_logic_vector(1 downto 0);
    signal ULT_u8_u1_101_wire : std_logic_vector(0 downto 0);
    signal ULT_u8_u1_108_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_95_data_0 : std_logic_vector(1 downto 0);
    signal array_obj_ref_95_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_95_index_partial_sum_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_95_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_95_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_95_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_95_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_95_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_95_word_offset_0 : std_logic_vector(3 downto 0);
    signal konst_100_wire_constant : std_logic_vector(7 downto 0);
    signal konst_107_wire_constant : std_logic_vector(7 downto 0);
    signal konst_77_wire_constant : std_logic_vector(7 downto 0);
    signal konst_90_wire_constant : std_logic_vector(7 downto 0);
    signal nI_79 : std_logic_vector(7 downto 0);
    signal nI_79_73_buffered : std_logic_vector(7 downto 0);
    signal nJ_92 : std_logic_vector(7 downto 0);
    signal nJ_92_86_buffered : std_logic_vector(7 downto 0);
    signal type_cast_72_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_85_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_ZERO_2_96_wire_constant <= "00";
    array_obj_ref_95_offset_scale_factor_0 <= "0100";
    array_obj_ref_95_offset_scale_factor_1 <= "0001";
    array_obj_ref_95_resized_base_address <= "0000";
    array_obj_ref_95_word_offset_0 <= "0000";
    konst_100_wire_constant <= "00000011";
    konst_107_wire_constant <= "00000011";
    konst_77_wire_constant <= "00000001";
    konst_90_wire_constant <= "00000001";
    type_cast_72_wire_constant <= "00000000";
    type_cast_85_wire_constant <= "00000000";
    phi_stmt_69: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_72_wire_constant & nI_79_73_buffered;
      req <= phi_stmt_69_req_0 & phi_stmt_69_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_69",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_69_ack_0,
          idata => idata,
          odata => I_69,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_69
    phi_stmt_82: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_85_wire_constant & nJ_92_86_buffered;
      req <= phi_stmt_82_req_0 & phi_stmt_82_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_82",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_82_ack_0,
          idata => idata,
          odata => J_82,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_82
    nI_79_73_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nI_79_73_buf_req_0;
      nI_79_73_buf_ack_0<= wack(0);
      rreq(0) <= nI_79_73_buf_req_1;
      nI_79_73_buf_ack_1<= rack(0);
      nI_79_73_buf : InterlockBuffer generic map ( -- 
        name => "nI_79_73_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nI_79,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nI_79_73_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nJ_92_86_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nJ_92_86_buf_req_0;
      nJ_92_86_buf_ack_0<= wack(0);
      rreq(0) <= nJ_92_86_buf_req_1;
      nJ_92_86_buf_ack_1<= rack(0);
      nJ_92_86_buf : InterlockBuffer generic map ( -- 
        name => "nJ_92_86_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nJ_92,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nJ_92_86_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_95_addr_0
    process(array_obj_ref_95_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_95_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_95_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_95_gather_scatter
    process(R_ZERO_2_96_wire_constant) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(1 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ZERO_2_96_wire_constant;
      ov(1 downto 0) := iv;
      array_obj_ref_95_data_0 <= ov(1 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_95_index_0_resize
    process(I_69) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_69;
      ov := iv(3 downto 0);
      R_I_93_resized <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_95_index_1_rename
    process(R_J_94_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_J_94_resized;
      ov(3 downto 0) := iv;
      R_J_94_scaled <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_95_index_1_resize
    process(J_82) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := J_82;
      ov := iv(3 downto 0);
      R_J_94_resized <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_95_index_offset
    process(array_obj_ref_95_index_partial_sum_1) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_95_index_partial_sum_1;
      ov(3 downto 0) := iv;
      array_obj_ref_95_final_offset <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_95_root_address_inst
    process(array_obj_ref_95_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_95_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_95_root_address <= ov(3 downto 0);
      --
    end process;
    if_stmt_105_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u8_u1_108_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_105_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_105_branch_req_0,
          ack0 => if_stmt_105_branch_ack_0,
          ack1 => if_stmt_105_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_98_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u8_u1_101_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_98_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_98_branch_req_0,
          ack0 => if_stmt_98_branch_ack_0,
          ack1 => if_stmt_98_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- flow through binary operator ADD_u8_u8_78_inst
    nI_79 <= std_logic_vector(unsigned(I_69) + unsigned(konst_77_wire_constant));
    -- flow through binary operator ADD_u8_u8_91_inst
    nJ_92 <= std_logic_vector(unsigned(J_82) + unsigned(konst_90_wire_constant));
    -- flow through binary operator ULT_u8_u1_101_inst
    process(J_82) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(J_82, konst_100_wire_constant, tmp_var);
      ULT_u8_u1_101_wire <= tmp_var; --
    end process;
    -- flow through binary operator ULT_u8_u1_108_inst
    process(I_69) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(I_69, konst_107_wire_constant, tmp_var);
      ULT_u8_u1_108_wire <= tmp_var; --
    end process;
    -- shared split operator group (4) : array_obj_ref_95_index_0_scale 
    ApIntMul_group_4: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_I_93_resized;
      R_I_93_scaled <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_95_index_0_scale_req_0;
      array_obj_ref_95_index_0_scale_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_95_index_0_scale_req_1;
      array_obj_ref_95_index_0_scale_ack_1 <= ackR_unguarded(0);
      ApIntMul_group_4_gI: SplitGuardInterface generic map(name => "ApIntMul_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          name => "ApIntMul_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0100",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : array_obj_ref_95_index_sum_1 
    ApIntAdd_group_5: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_J_94_scaled & R_I_93_scaled;
      array_obj_ref_95_index_partial_sum_1 <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_95_index_sum_1_req_0;
      array_obj_ref_95_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_95_index_sum_1_req_1;
      array_obj_ref_95_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_5_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_5",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 4, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared store operator group (0) : array_obj_ref_95_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(3 downto 0);
      signal data_in: std_logic_vector(1 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_95_store_0_req_0;
      array_obj_ref_95_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_95_store_0_req_1;
      array_obj_ref_95_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_95_word_address_0;
      data_in <= array_obj_ref_95_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 4,
        data_width => 2,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(3 downto 0),
          mdata => memory_space_0_sr_data(1 downto 0),
          mtag => memory_space_0_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end initialiseCounters_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity inputPort_1_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    in_data_1_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_1_pipe_read_data : in   std_logic_vector(31 downto 0);
    noblock_obuf_1_3_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_3_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_1_4_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_4_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_1_1_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_1_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_1_2_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_2_pipe_write_data : out  std_logic_vector(32 downto 0);
    updateCounter_call_reqs : out  std_logic_vector(0 downto 0);
    updateCounter_call_acks : in   std_logic_vector(0 downto 0);
    updateCounter_call_data : out  std_logic_vector(16 downto 0);
    updateCounter_call_tag  :  out  std_logic_vector(0 downto 0);
    updateCounter_return_reqs : out  std_logic_vector(0 downto 0);
    updateCounter_return_acks : in   std_logic_vector(0 downto 0);
    updateCounter_return_data : in   std_logic_vector(0 downto 0);
    updateCounter_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity inputPort_1_Daemon;
architecture inputPort_1_Daemon_arch of inputPort_1_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal inputPort_1_Daemon_CP_1105_start: Boolean;
  signal inputPort_1_Daemon_CP_1105_symbol: Boolean;
  -- volatile/operator module components. 
  component updateCounter is -- 
    generic (tag_length : integer); 
    port ( -- 
      input_port : in  std_logic_vector(7 downto 0);
      output_port : in  std_logic_vector(7 downto 0);
      up : in  std_logic_vector(0 downto 0);
      continue : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(3 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(1 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(1 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal RPIPE_in_data_1_223_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_1_2_334_inst_ack_0 : boolean;
  signal EQ_u8_u1_296_inst_ack_1 : boolean;
  signal RPIPE_in_data_1_223_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_1_1_327_inst_ack_1 : boolean;
  signal EQ_u8_u1_296_inst_req_0 : boolean;
  signal do_while_stmt_215_branch_req_0 : boolean;
  signal phi_stmt_217_req_1 : boolean;
  signal EQ_u8_u1_296_inst_req_1 : boolean;
  signal phi_stmt_224_req_0 : boolean;
  signal WPIPE_noblock_obuf_1_2_334_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_1_1_327_inst_req_1 : boolean;
  signal RPIPE_in_data_1_223_inst_ack_0 : boolean;
  signal phi_stmt_224_req_1 : boolean;
  signal W_data_to_outport_317_delayed_4_0_330_inst_ack_0 : boolean;
  signal RPIPE_in_data_1_223_inst_req_1 : boolean;
  signal W_data_to_outport_317_delayed_4_0_330_inst_req_1 : boolean;
  signal W_data_to_outport_317_delayed_4_0_330_inst_ack_1 : boolean;
  signal EQ_u8_u1_296_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_1_1_327_inst_ack_0 : boolean;
  signal W_data_to_outport_313_delayed_4_0_323_inst_ack_0 : boolean;
  signal W_data_to_outport_317_delayed_4_0_330_inst_req_0 : boolean;
  signal EQ_u8_u1_286_inst_ack_1 : boolean;
  signal phi_stmt_224_ack_0 : boolean;
  signal phi_stmt_217_ack_0 : boolean;
  signal WPIPE_noblock_obuf_1_1_327_inst_req_0 : boolean;
  signal phi_stmt_217_req_0 : boolean;
  signal W_data_to_outport_313_delayed_4_0_323_inst_ack_1 : boolean;
  signal EQ_u8_u1_306_inst_req_1 : boolean;
  signal next_last_dest_id_268_226_buf_req_0 : boolean;
  signal next_last_dest_id_268_226_buf_ack_0 : boolean;
  signal EQ_u8_u1_316_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_1_2_334_inst_ack_1 : boolean;
  signal next_last_dest_id_268_226_buf_req_1 : boolean;
  signal next_last_dest_id_268_226_buf_ack_1 : boolean;
  signal EQ_u8_u1_306_inst_ack_1 : boolean;
  signal W_data_to_outport_313_delayed_4_0_323_inst_req_0 : boolean;
  signal EQ_u8_u1_316_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_1_2_334_inst_req_1 : boolean;
  signal EQ_u8_u1_316_inst_req_0 : boolean;
  signal call_updateCounter_expr_281_inst_req_0 : boolean;
  signal call_updateCounter_expr_281_inst_ack_0 : boolean;
  signal next_count_down_262_219_buf_req_0 : boolean;
  signal call_updateCounter_expr_281_inst_req_1 : boolean;
  signal call_updateCounter_expr_281_inst_ack_1 : boolean;
  signal EQ_u8_u1_306_inst_req_0 : boolean;
  signal next_count_down_262_219_buf_ack_0 : boolean;
  signal next_count_down_262_219_buf_req_1 : boolean;
  signal next_count_down_262_219_buf_ack_1 : boolean;
  signal EQ_u8_u1_286_inst_req_0 : boolean;
  signal EQ_u8_u1_306_inst_ack_0 : boolean;
  signal EQ_u8_u1_286_inst_ack_0 : boolean;
  signal EQ_u8_u1_316_inst_ack_0 : boolean;
  signal W_data_to_outport_313_delayed_4_0_323_inst_req_1 : boolean;
  signal EQ_u8_u1_286_inst_req_1 : boolean;
  signal W_data_to_outport_321_delayed_4_0_337_inst_req_0 : boolean;
  signal W_data_to_outport_321_delayed_4_0_337_inst_ack_0 : boolean;
  signal W_data_to_outport_321_delayed_4_0_337_inst_req_1 : boolean;
  signal W_data_to_outport_321_delayed_4_0_337_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_1_3_341_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_1_3_341_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_1_3_341_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_1_3_341_inst_ack_1 : boolean;
  signal W_data_to_outport_325_delayed_4_0_344_inst_req_0 : boolean;
  signal W_data_to_outport_325_delayed_4_0_344_inst_ack_0 : boolean;
  signal W_data_to_outport_325_delayed_4_0_344_inst_req_1 : boolean;
  signal W_data_to_outport_325_delayed_4_0_344_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_1_4_348_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_1_4_348_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_1_4_348_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_1_4_348_inst_ack_1 : boolean;
  signal do_while_stmt_215_branch_ack_0 : boolean;
  signal do_while_stmt_215_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "inputPort_1_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  inputPort_1_Daemon_CP_1105_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "inputPort_1_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_1_Daemon_CP_1105_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= inputPort_1_Daemon_CP_1105_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_1_Daemon_CP_1105_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  inputPort_1_Daemon_CP_1105: Block -- control-path 
    signal inputPort_1_Daemon_CP_1105_elements: BooleanArray(105 downto 0);
    -- 
  begin -- 
    inputPort_1_Daemon_CP_1105_elements(0) <= inputPort_1_Daemon_CP_1105_start;
    inputPort_1_Daemon_CP_1105_symbol <= inputPort_1_Daemon_CP_1105_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_214/$entry
      -- CP-element group 0: 	 branch_block_stmt_214/branch_block_stmt_214__entry__
      -- CP-element group 0: 	 branch_block_stmt_214/do_while_stmt_215__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	105 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_214/$exit
      -- CP-element group 1: 	 branch_block_stmt_214/branch_block_stmt_214__exit__
      -- CP-element group 1: 	 branch_block_stmt_214/do_while_stmt_215__exit__
      -- 
    inputPort_1_Daemon_CP_1105_elements(1) <= inputPort_1_Daemon_CP_1105_elements(105);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_214/do_while_stmt_215/$entry
      -- CP-element group 2: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215__entry__
      -- 
    inputPort_1_Daemon_CP_1105_elements(2) <= inputPort_1_Daemon_CP_1105_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	105 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215__exit__
      -- 
    -- Element group inputPort_1_Daemon_CP_1105_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_214/do_while_stmt_215/loop_back
      -- 
    -- Element group inputPort_1_Daemon_CP_1105_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	103 
    -- CP-element group 5: 	104 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_214/do_while_stmt_215/condition_done
      -- CP-element group 5: 	 branch_block_stmt_214/do_while_stmt_215/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_214/do_while_stmt_215/loop_taken/$entry
      -- 
    inputPort_1_Daemon_CP_1105_elements(5) <= inputPort_1_Daemon_CP_1105_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	102 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_214/do_while_stmt_215/loop_body_done
      -- 
    inputPort_1_Daemon_CP_1105_elements(6) <= inputPort_1_Daemon_CP_1105_elements(102);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	21 
    -- CP-element group 7: 	44 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/back_edge_to_loop_body
      -- 
    inputPort_1_Daemon_CP_1105_elements(7) <= inputPort_1_Daemon_CP_1105_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	23 
    -- CP-element group 8: 	46 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/first_time_through_loop_body
      -- 
    inputPort_1_Daemon_CP_1105_elements(8) <= inputPort_1_Daemon_CP_1105_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	39 
    -- CP-element group 9: 	40 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	17 
    -- CP-element group 9: 	101 
    -- CP-element group 9: 	34 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_221_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/$entry
      -- 
    -- Element group inputPort_1_Daemon_CP_1105_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	101 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/condition_evaluated
      -- 
    condition_evaluated_1129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(10), ack => do_while_stmt_215_branch_req_0); -- 
    inputPort_1_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_1105_elements(15) & inputPort_1_Daemon_CP_1105_elements(101);
      gj_inputPort_1_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	39 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	16 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	18 
    -- CP-element group 11: 	35 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_224_sample_start__ps
      -- CP-element group 11: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/aggregated_phi_sample_req
      -- 
    inputPort_1_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 7,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_1105_elements(39) & inputPort_1_Daemon_CP_1105_elements(9) & inputPort_1_Daemon_CP_1105_elements(16) & inputPort_1_Daemon_CP_1105_elements(15);
      gj_inputPort_1_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	37 
    -- CP-element group 12: 	19 
    -- CP-element group 12: 	41 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12: 	102 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	39 
    -- CP-element group 12: 	16 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_221_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_224_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_217_sample_completed_
      -- 
    inputPort_1_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_1105_elements(37) & inputPort_1_Daemon_CP_1105_elements(19) & inputPort_1_Daemon_CP_1105_elements(41);
      gj_inputPort_1_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	102 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/aggregated_phi_sample_ack_d
      -- 
    -- Element group inputPort_1_Daemon_CP_1105_elements(13) is a control-delay.
    cp_element_13_delay: control_delay_element  generic map(name => " 13_delay", delay_value => 1)  port map(req => inputPort_1_Daemon_CP_1105_elements(12), ack => inputPort_1_Daemon_CP_1105_elements(13), clk => clk, reset =>reset);
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	40 
    -- CP-element group 14: 	17 
    -- CP-element group 14: 	34 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	42 
    -- CP-element group 14: 	36 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_217_update_start__ps
      -- CP-element group 14: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/aggregated_phi_update_req
      -- 
    inputPort_1_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_1105_elements(40) & inputPort_1_Daemon_CP_1105_elements(17) & inputPort_1_Daemon_CP_1105_elements(34);
      gj_inputPort_1_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	38 
    -- CP-element group 15: 	20 
    -- CP-element group 15: 	43 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/aggregated_phi_update_ack
      -- 
    inputPort_1_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_1105_elements(38) & inputPort_1_Daemon_CP_1105_elements(20) & inputPort_1_Daemon_CP_1105_elements(43);
      gj_inputPort_1_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	11 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_217_sample_start_
      -- 
    inputPort_1_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_1105_elements(9) & inputPort_1_Daemon_CP_1105_elements(12);
      gj_inputPort_1_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	9 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	59 
    -- CP-element group 17: 	63 
    -- CP-element group 17: 	67 
    -- CP-element group 17: 	71 
    -- CP-element group 17: 	75 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	14 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_217_update_start_
      -- 
    inputPort_1_Daemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_1105_elements(9) & inputPort_1_Daemon_CP_1105_elements(59) & inputPort_1_Daemon_CP_1105_elements(63) & inputPort_1_Daemon_CP_1105_elements(67) & inputPort_1_Daemon_CP_1105_elements(71) & inputPort_1_Daemon_CP_1105_elements(75);
      gj_inputPort_1_Daemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	11 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_217_sample_start__ps
      -- 
    inputPort_1_Daemon_CP_1105_elements(18) <= inputPort_1_Daemon_CP_1105_elements(11);
    -- CP-element group 19:  join  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	12 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_217_sample_completed__ps
      -- 
    -- Element group inputPort_1_Daemon_CP_1105_elements(19) is bound as output of CP function.
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: 	57 
    -- CP-element group 20: 	61 
    -- CP-element group 20: 	65 
    -- CP-element group 20: 	69 
    -- CP-element group 20: 	73 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_217_update_completed__ps
      -- CP-element group 20: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_217_update_completed_
      -- 
    -- Element group inputPort_1_Daemon_CP_1105_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	7 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_217_loopback_trigger
      -- 
    inputPort_1_Daemon_CP_1105_elements(21) <= inputPort_1_Daemon_CP_1105_elements(7);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_217_loopback_sample_req
      -- CP-element group 22: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_217_loopback_sample_req_ps
      -- 
    phi_stmt_217_loopback_sample_req_1145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_217_loopback_sample_req_1145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(22), ack => phi_stmt_217_req_0); -- 
    -- Element group inputPort_1_Daemon_CP_1105_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	8 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_217_entry_trigger
      -- 
    inputPort_1_Daemon_CP_1105_elements(23) <= inputPort_1_Daemon_CP_1105_elements(8);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_217_entry_sample_req
      -- CP-element group 24: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_217_entry_sample_req_ps
      -- 
    phi_stmt_217_entry_sample_req_1148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_217_entry_sample_req_1148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(24), ack => phi_stmt_217_req_1); -- 
    -- Element group inputPort_1_Daemon_CP_1105_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_217_phi_mux_ack_ps
      -- CP-element group 25: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_217_phi_mux_ack
      -- 
    phi_stmt_217_phi_mux_ack_1151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_217_ack_0, ack => inputPort_1_Daemon_CP_1105_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_count_down_219_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_count_down_219_sample_start__ps
      -- CP-element group 26: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_count_down_219_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_count_down_219_Sample/req
      -- 
    req_1164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(26), ack => next_count_down_262_219_buf_req_0); -- 
    -- Element group inputPort_1_Daemon_CP_1105_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_count_down_219_update_start__ps
      -- CP-element group 27: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_count_down_219_update_start_
      -- CP-element group 27: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_count_down_219_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_count_down_219_Update/req
      -- 
    req_1169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(27), ack => next_count_down_262_219_buf_req_1); -- 
    -- Element group inputPort_1_Daemon_CP_1105_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_count_down_219_sample_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_count_down_219_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_count_down_219_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_count_down_219_Sample/ack
      -- 
    ack_1165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_262_219_buf_ack_0, ack => inputPort_1_Daemon_CP_1105_elements(28)); -- 
    -- CP-element group 29:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_count_down_219_update_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_count_down_219_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_count_down_219_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_count_down_219_Update/ack
      -- 
    ack_1170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_262_219_buf_ack_1, ack => inputPort_1_Daemon_CP_1105_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_ZERO_16_220_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_ZERO_16_220_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_ZERO_16_220_sample_start__ps
      -- CP-element group 30: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_ZERO_16_220_sample_completed__ps
      -- 
    -- Element group inputPort_1_Daemon_CP_1105_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_ZERO_16_220_update_start_
      -- CP-element group 31: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_ZERO_16_220_update_start__ps
      -- 
    -- Element group inputPort_1_Daemon_CP_1105_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	33 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_ZERO_16_220_update_completed__ps
      -- 
    inputPort_1_Daemon_CP_1105_elements(32) <= inputPort_1_Daemon_CP_1105_elements(33);
    -- CP-element group 33:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	32 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_ZERO_16_220_update_completed_
      -- 
    -- Element group inputPort_1_Daemon_CP_1105_elements(33) is a control-delay.
    cp_element_33_delay: control_delay_element  generic map(name => " 33_delay", delay_value => 1)  port map(req => inputPort_1_Daemon_CP_1105_elements(31), ack => inputPort_1_Daemon_CP_1105_elements(33), clk => clk, reset =>reset);
    -- CP-element group 34:  join  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	9 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	59 
    -- CP-element group 34: 	90 
    -- CP-element group 34: 	96 
    -- CP-element group 34: 	63 
    -- CP-element group 34: 	67 
    -- CP-element group 34: 	71 
    -- CP-element group 34: 	75 
    -- CP-element group 34: 	78 
    -- CP-element group 34: 	84 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	14 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_221_update_start_
      -- 
    inputPort_1_Daemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_1105_elements(9) & inputPort_1_Daemon_CP_1105_elements(59) & inputPort_1_Daemon_CP_1105_elements(90) & inputPort_1_Daemon_CP_1105_elements(96) & inputPort_1_Daemon_CP_1105_elements(63) & inputPort_1_Daemon_CP_1105_elements(67) & inputPort_1_Daemon_CP_1105_elements(71) & inputPort_1_Daemon_CP_1105_elements(75) & inputPort_1_Daemon_CP_1105_elements(78) & inputPort_1_Daemon_CP_1105_elements(84);
      gj_inputPort_1_Daemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	11 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	38 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/RPIPE_in_data_1_223_Sample/rr
      -- CP-element group 35: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/RPIPE_in_data_1_223_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/RPIPE_in_data_1_223_sample_start_
      -- 
    rr_1191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(35), ack => RPIPE_in_data_1_223_inst_req_0); -- 
    inputPort_1_Daemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_1105_elements(11) & inputPort_1_Daemon_CP_1105_elements(38);
      gj_inputPort_1_Daemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	37 
    -- CP-element group 36: 	14 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/RPIPE_in_data_1_223_Update/cr
      -- CP-element group 36: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/RPIPE_in_data_1_223_update_start_
      -- CP-element group 36: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/RPIPE_in_data_1_223_Update/$entry
      -- 
    cr_1196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(36), ack => RPIPE_in_data_1_223_inst_req_1); -- 
    inputPort_1_Daemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_1105_elements(37) & inputPort_1_Daemon_CP_1105_elements(14);
      gj_inputPort_1_Daemon_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	12 
    -- CP-element group 37: 	36 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/RPIPE_in_data_1_223_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/RPIPE_in_data_1_223_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/RPIPE_in_data_1_223_sample_completed_
      -- 
    ra_1192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_1_223_inst_ack_0, ack => inputPort_1_Daemon_CP_1105_elements(37)); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	15 
    -- CP-element group 38: 	57 
    -- CP-element group 38: 	90 
    -- CP-element group 38: 	96 
    -- CP-element group 38: 	61 
    -- CP-element group 38: 	65 
    -- CP-element group 38: 	69 
    -- CP-element group 38: 	73 
    -- CP-element group 38: 	78 
    -- CP-element group 38: 	84 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	35 
    -- CP-element group 38:  members (16) 
      -- CP-element group 38: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/RPIPE_in_data_1_223_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_325_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_332_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_332_Sample/req
      -- CP-element group 38: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/RPIPE_in_data_1_223_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/RPIPE_in_data_1_223_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_325_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_325_Sample/req
      -- CP-element group 38: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_221_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_332_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_339_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_339_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_339_Sample/req
      -- CP-element group 38: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_346_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_346_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_346_Sample/req
      -- 
    ca_1197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_1_223_inst_ack_1, ack => inputPort_1_Daemon_CP_1105_elements(38)); -- 
    req_1375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(38), ack => W_data_to_outport_321_delayed_4_0_337_inst_req_0); -- 
    req_1403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(38), ack => W_data_to_outport_325_delayed_4_0_344_inst_req_0); -- 
    req_1319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(38), ack => W_data_to_outport_313_delayed_4_0_323_inst_req_0); -- 
    req_1347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(38), ack => W_data_to_outport_317_delayed_4_0_330_inst_req_0); -- 
    -- CP-element group 39:  join  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	9 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	12 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	11 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_224_sample_start_
      -- 
    inputPort_1_Daemon_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_1105_elements(9) & inputPort_1_Daemon_CP_1105_elements(12);
      gj_inputPort_1_Daemon_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	9 
    -- CP-element group 40: marked-predecessors 
    -- CP-element group 40: 	59 
    -- CP-element group 40: 	63 
    -- CP-element group 40: 	67 
    -- CP-element group 40: 	71 
    -- CP-element group 40: 	75 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	14 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_224_update_start_
      -- 
    inputPort_1_Daemon_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_1105_elements(9) & inputPort_1_Daemon_CP_1105_elements(59) & inputPort_1_Daemon_CP_1105_elements(63) & inputPort_1_Daemon_CP_1105_elements(67) & inputPort_1_Daemon_CP_1105_elements(71) & inputPort_1_Daemon_CP_1105_elements(75);
      gj_inputPort_1_Daemon_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	12 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_224_sample_completed__ps
      -- 
    -- Element group inputPort_1_Daemon_CP_1105_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	14 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_224_update_start__ps
      -- 
    inputPort_1_Daemon_CP_1105_elements(42) <= inputPort_1_Daemon_CP_1105_elements(14);
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	15 
    -- CP-element group 43: 	57 
    -- CP-element group 43: 	61 
    -- CP-element group 43: 	65 
    -- CP-element group 43: 	69 
    -- CP-element group 43: 	73 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_224_update_completed__ps
      -- CP-element group 43: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_224_update_completed_
      -- 
    -- Element group inputPort_1_Daemon_CP_1105_elements(43) is bound as output of CP function.
    -- CP-element group 44:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	7 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_224_loopback_trigger
      -- 
    inputPort_1_Daemon_CP_1105_elements(44) <= inputPort_1_Daemon_CP_1105_elements(7);
    -- CP-element group 45:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_224_loopback_sample_req
      -- CP-element group 45: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_224_loopback_sample_req_ps
      -- 
    phi_stmt_224_loopback_sample_req_1207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_224_loopback_sample_req_1207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(45), ack => phi_stmt_224_req_0); -- 
    -- Element group inputPort_1_Daemon_CP_1105_elements(45) is bound as output of CP function.
    -- CP-element group 46:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	8 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_224_entry_trigger
      -- 
    inputPort_1_Daemon_CP_1105_elements(46) <= inputPort_1_Daemon_CP_1105_elements(8);
    -- CP-element group 47:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_224_entry_sample_req
      -- CP-element group 47: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_224_entry_sample_req_ps
      -- 
    phi_stmt_224_entry_sample_req_1210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_224_entry_sample_req_1210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(47), ack => phi_stmt_224_req_1); -- 
    -- Element group inputPort_1_Daemon_CP_1105_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_224_phi_mux_ack
      -- CP-element group 48: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/phi_stmt_224_phi_mux_ack_ps
      -- 
    phi_stmt_224_phi_mux_ack_1213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_224_ack_0, ack => inputPort_1_Daemon_CP_1105_elements(48)); -- 
    -- CP-element group 49:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_last_dest_id_226_sample_start__ps
      -- CP-element group 49: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_last_dest_id_226_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_last_dest_id_226_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_last_dest_id_226_Sample/req
      -- 
    req_1226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(49), ack => next_last_dest_id_268_226_buf_req_0); -- 
    -- Element group inputPort_1_Daemon_CP_1105_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_last_dest_id_226_update_start__ps
      -- CP-element group 50: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_last_dest_id_226_update_start_
      -- CP-element group 50: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_last_dest_id_226_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_last_dest_id_226_Update/req
      -- 
    req_1231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(50), ack => next_last_dest_id_268_226_buf_req_1); -- 
    -- Element group inputPort_1_Daemon_CP_1105_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_last_dest_id_226_sample_completed__ps
      -- CP-element group 51: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_last_dest_id_226_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_last_dest_id_226_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_last_dest_id_226_Sample/ack
      -- 
    ack_1227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_268_226_buf_ack_0, ack => inputPort_1_Daemon_CP_1105_elements(51)); -- 
    -- CP-element group 52:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_last_dest_id_226_update_completed__ps
      -- CP-element group 52: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_last_dest_id_226_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_last_dest_id_226_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/R_next_last_dest_id_226_Update/ack
      -- 
    ack_1232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_268_226_buf_ack_1, ack => inputPort_1_Daemon_CP_1105_elements(52)); -- 
    -- CP-element group 53:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/konst_227_sample_start__ps
      -- CP-element group 53: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/konst_227_sample_completed__ps
      -- CP-element group 53: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/konst_227_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/konst_227_sample_completed_
      -- 
    -- Element group inputPort_1_Daemon_CP_1105_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (2) 
      -- CP-element group 54: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/konst_227_update_start__ps
      -- CP-element group 54: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/konst_227_update_start_
      -- 
    -- Element group inputPort_1_Daemon_CP_1105_elements(54) is bound as output of CP function.
    -- CP-element group 55:  join  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/konst_227_update_completed__ps
      -- 
    inputPort_1_Daemon_CP_1105_elements(55) <= inputPort_1_Daemon_CP_1105_elements(56);
    -- CP-element group 56:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	55 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/konst_227_update_completed_
      -- 
    -- Element group inputPort_1_Daemon_CP_1105_elements(56) is a control-delay.
    cp_element_56_delay: control_delay_element  generic map(name => " 56_delay", delay_value => 1)  port map(req => inputPort_1_Daemon_CP_1105_elements(54), ack => inputPort_1_Daemon_CP_1105_elements(56), clk => clk, reset =>reset);
    -- CP-element group 57:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	38 
    -- CP-element group 57: 	20 
    -- CP-element group 57: 	43 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/call_updateCounter_expr_281_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/call_updateCounter_expr_281_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/call_updateCounter_expr_281_Sample/req
      -- 
    req_1249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(57), ack => call_updateCounter_expr_281_inst_req_0); -- 
    inputPort_1_Daemon_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_1105_elements(38) & inputPort_1_Daemon_CP_1105_elements(20) & inputPort_1_Daemon_CP_1105_elements(43);
      gj_inputPort_1_Daemon_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	87 
    -- CP-element group 58: 	93 
    -- CP-element group 58: 	99 
    -- CP-element group 58: 	81 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/call_updateCounter_expr_281_update_start_
      -- CP-element group 58: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/call_updateCounter_expr_281_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/call_updateCounter_expr_281_Update/req
      -- 
    req_1254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(58), ack => call_updateCounter_expr_281_inst_req_1); -- 
    inputPort_1_Daemon_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_1105_elements(87) & inputPort_1_Daemon_CP_1105_elements(93) & inputPort_1_Daemon_CP_1105_elements(99) & inputPort_1_Daemon_CP_1105_elements(81);
      gj_inputPort_1_Daemon_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: marked-successors 
    -- CP-element group 59: 	40 
    -- CP-element group 59: 	17 
    -- CP-element group 59: 	34 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/call_updateCounter_expr_281_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/call_updateCounter_expr_281_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/call_updateCounter_expr_281_Sample/ack
      -- 
    ack_1250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_updateCounter_expr_281_inst_ack_0, ack => inputPort_1_Daemon_CP_1105_elements(59)); -- 
    -- CP-element group 60:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	92 
    -- CP-element group 60: 	98 
    -- CP-element group 60: 	80 
    -- CP-element group 60: 	86 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/call_updateCounter_expr_281_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/call_updateCounter_expr_281_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/call_updateCounter_expr_281_Update/ack
      -- 
    ack_1255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_updateCounter_expr_281_inst_ack_1, ack => inputPort_1_Daemon_CP_1105_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	38 
    -- CP-element group 61: 	20 
    -- CP-element group 61: 	43 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_286_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_286_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_286_Sample/rr
      -- 
    rr_1263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(61), ack => EQ_u8_u1_286_inst_req_0); -- 
    inputPort_1_Daemon_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_1105_elements(38) & inputPort_1_Daemon_CP_1105_elements(20) & inputPort_1_Daemon_CP_1105_elements(43);
      gj_inputPort_1_Daemon_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	81 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_286_update_start_
      -- CP-element group 62: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_286_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_286_Update/cr
      -- 
    cr_1268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(62), ack => EQ_u8_u1_286_inst_req_1); -- 
    inputPort_1_Daemon_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_1_Daemon_CP_1105_elements(81);
      gj_inputPort_1_Daemon_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	40 
    -- CP-element group 63: 	17 
    -- CP-element group 63: 	34 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_286_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_286_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_286_Sample/ra
      -- 
    ra_1264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_286_inst_ack_0, ack => inputPort_1_Daemon_CP_1105_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	80 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_286_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_286_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_286_Update/$exit
      -- 
    ca_1269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_286_inst_ack_1, ack => inputPort_1_Daemon_CP_1105_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	38 
    -- CP-element group 65: 	20 
    -- CP-element group 65: 	43 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_296_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_296_Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_296_Sample/$entry
      -- 
    rr_1277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(65), ack => EQ_u8_u1_296_inst_req_0); -- 
    inputPort_1_Daemon_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_1105_elements(38) & inputPort_1_Daemon_CP_1105_elements(20) & inputPort_1_Daemon_CP_1105_elements(43);
      gj_inputPort_1_Daemon_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	87 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_296_Update/cr
      -- CP-element group 66: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_296_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_296_update_start_
      -- 
    cr_1282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(66), ack => EQ_u8_u1_296_inst_req_1); -- 
    inputPort_1_Daemon_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_1_Daemon_CP_1105_elements(87);
      gj_inputPort_1_Daemon_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	40 
    -- CP-element group 67: 	17 
    -- CP-element group 67: 	34 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_296_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_296_Sample/ra
      -- CP-element group 67: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_296_Sample/$exit
      -- 
    ra_1278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_296_inst_ack_0, ack => inputPort_1_Daemon_CP_1105_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	86 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_296_Update/ca
      -- CP-element group 68: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_296_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_296_Update/$exit
      -- 
    ca_1283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_296_inst_ack_1, ack => inputPort_1_Daemon_CP_1105_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	38 
    -- CP-element group 69: 	20 
    -- CP-element group 69: 	43 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_306_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_306_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_306_Sample/rr
      -- 
    rr_1291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(69), ack => EQ_u8_u1_306_inst_req_0); -- 
    inputPort_1_Daemon_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_1105_elements(38) & inputPort_1_Daemon_CP_1105_elements(20) & inputPort_1_Daemon_CP_1105_elements(43);
      gj_inputPort_1_Daemon_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	93 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_306_update_start_
      -- CP-element group 70: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_306_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_306_Update/$entry
      -- 
    cr_1296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(70), ack => EQ_u8_u1_306_inst_req_1); -- 
    inputPort_1_Daemon_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_1_Daemon_CP_1105_elements(93);
      gj_inputPort_1_Daemon_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: marked-successors 
    -- CP-element group 71: 	40 
    -- CP-element group 71: 	17 
    -- CP-element group 71: 	34 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_306_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_306_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_306_Sample/ra
      -- 
    ra_1292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_306_inst_ack_0, ack => inputPort_1_Daemon_CP_1105_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	92 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_306_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_306_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_306_Update/ca
      -- 
    ca_1297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_306_inst_ack_1, ack => inputPort_1_Daemon_CP_1105_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	38 
    -- CP-element group 73: 	20 
    -- CP-element group 73: 	43 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_316_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_316_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_316_Sample/rr
      -- 
    rr_1305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(73), ack => EQ_u8_u1_316_inst_req_0); -- 
    inputPort_1_Daemon_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_1105_elements(38) & inputPort_1_Daemon_CP_1105_elements(20) & inputPort_1_Daemon_CP_1105_elements(43);
      gj_inputPort_1_Daemon_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	99 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_316_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_316_update_start_
      -- CP-element group 74: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_316_Update/cr
      -- 
    cr_1310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(74), ack => EQ_u8_u1_316_inst_req_1); -- 
    inputPort_1_Daemon_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_1_Daemon_CP_1105_elements(99);
      gj_inputPort_1_Daemon_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	40 
    -- CP-element group 75: 	17 
    -- CP-element group 75: 	34 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_316_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_316_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_316_Sample/ra
      -- 
    ra_1306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_316_inst_ack_0, ack => inputPort_1_Daemon_CP_1105_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	98 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_316_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_316_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/EQ_u8_u1_316_Update/ca
      -- 
    ca_1311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_316_inst_ack_1, ack => inputPort_1_Daemon_CP_1105_elements(76)); -- 
    -- CP-element group 77:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	81 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_325_update_start_
      -- CP-element group 77: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_325_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_325_Update/req
      -- 
    req_1324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(77), ack => W_data_to_outport_313_delayed_4_0_323_inst_req_1); -- 
    inputPort_1_Daemon_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_1_Daemon_CP_1105_elements(81);
      gj_inputPort_1_Daemon_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	38 
    -- CP-element group 78: successors 
    -- CP-element group 78: marked-successors 
    -- CP-element group 78: 	34 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_325_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_325_Sample/ack
      -- CP-element group 78: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_325_Sample/$exit
      -- 
    ack_1320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_313_delayed_4_0_323_inst_ack_0, ack => inputPort_1_Daemon_CP_1105_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_325_Update/ack
      -- CP-element group 79: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_325_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_325_Update/$exit
      -- 
    ack_1325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_313_delayed_4_0_323_inst_ack_1, ack => inputPort_1_Daemon_CP_1105_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	60 
    -- CP-element group 80: 	64 
    -- CP-element group 80: 	79 
    -- CP-element group 80: marked-predecessors 
    -- CP-element group 80: 	82 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_1_327_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_1_327_Sample/req
      -- CP-element group 80: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_1_327_sample_start_
      -- 
    req_1333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(80), ack => WPIPE_noblock_obuf_1_1_327_inst_req_0); -- 
    inputPort_1_Daemon_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_1105_elements(60) & inputPort_1_Daemon_CP_1105_elements(64) & inputPort_1_Daemon_CP_1105_elements(79) & inputPort_1_Daemon_CP_1105_elements(82);
      gj_inputPort_1_Daemon_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81: marked-successors 
    -- CP-element group 81: 	58 
    -- CP-element group 81: 	62 
    -- CP-element group 81: 	77 
    -- CP-element group 81:  members (6) 
      -- CP-element group 81: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_1_327_Update/req
      -- CP-element group 81: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_1_327_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_1_327_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_1_327_Sample/ack
      -- CP-element group 81: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_1_327_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_1_327_update_start_
      -- 
    ack_1334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_1_327_inst_ack_0, ack => inputPort_1_Daemon_CP_1105_elements(81)); -- 
    req_1338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(81), ack => WPIPE_noblock_obuf_1_1_327_inst_req_1); -- 
    -- CP-element group 82:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	102 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	80 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_1_327_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_1_327_Update/ack
      -- CP-element group 82: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_1_327_update_completed_
      -- 
    ack_1339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_1_327_inst_ack_1, ack => inputPort_1_Daemon_CP_1105_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: marked-predecessors 
    -- CP-element group 83: 	87 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_332_Update/req
      -- CP-element group 83: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_332_update_start_
      -- CP-element group 83: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_332_Update/$entry
      -- 
    req_1352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(83), ack => W_data_to_outport_317_delayed_4_0_330_inst_req_1); -- 
    inputPort_1_Daemon_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_1_Daemon_CP_1105_elements(87);
      gj_inputPort_1_Daemon_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	38 
    -- CP-element group 84: successors 
    -- CP-element group 84: marked-successors 
    -- CP-element group 84: 	34 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_332_Sample/ack
      -- CP-element group 84: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_332_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_332_sample_completed_
      -- 
    ack_1348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_317_delayed_4_0_330_inst_ack_0, ack => inputPort_1_Daemon_CP_1105_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_332_Update/ack
      -- CP-element group 85: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_332_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_332_Update/$exit
      -- 
    ack_1353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_317_delayed_4_0_330_inst_ack_1, ack => inputPort_1_Daemon_CP_1105_elements(85)); -- 
    -- CP-element group 86:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	60 
    -- CP-element group 86: 	68 
    -- CP-element group 86: 	85 
    -- CP-element group 86: marked-predecessors 
    -- CP-element group 86: 	88 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_2_334_Sample/req
      -- CP-element group 86: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_2_334_Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_2_334_sample_start_
      -- 
    req_1361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(86), ack => WPIPE_noblock_obuf_1_2_334_inst_req_0); -- 
    inputPort_1_Daemon_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_1105_elements(60) & inputPort_1_Daemon_CP_1105_elements(68) & inputPort_1_Daemon_CP_1105_elements(85) & inputPort_1_Daemon_CP_1105_elements(88);
      gj_inputPort_1_Daemon_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: marked-successors 
    -- CP-element group 87: 	58 
    -- CP-element group 87: 	66 
    -- CP-element group 87: 	83 
    -- CP-element group 87:  members (6) 
      -- CP-element group 87: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_2_334_Sample/ack
      -- CP-element group 87: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_2_334_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_2_334_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_2_334_update_start_
      -- CP-element group 87: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_2_334_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_2_334_Update/req
      -- 
    ack_1362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_2_334_inst_ack_0, ack => inputPort_1_Daemon_CP_1105_elements(87)); -- 
    req_1366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(87), ack => WPIPE_noblock_obuf_1_2_334_inst_req_1); -- 
    -- CP-element group 88:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	102 
    -- CP-element group 88: marked-successors 
    -- CP-element group 88: 	86 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_2_334_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_2_334_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_2_334_Update/ack
      -- 
    ack_1367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_2_334_inst_ack_1, ack => inputPort_1_Daemon_CP_1105_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	93 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_339_update_start_
      -- CP-element group 89: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_339_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_339_Update/req
      -- 
    req_1380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(89), ack => W_data_to_outport_321_delayed_4_0_337_inst_req_1); -- 
    inputPort_1_Daemon_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_1_Daemon_CP_1105_elements(93);
      gj_inputPort_1_Daemon_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	38 
    -- CP-element group 90: successors 
    -- CP-element group 90: marked-successors 
    -- CP-element group 90: 	34 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_339_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_339_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_339_Sample/ack
      -- 
    ack_1376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_321_delayed_4_0_337_inst_ack_0, ack => inputPort_1_Daemon_CP_1105_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_339_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_339_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_339_Update/ack
      -- 
    ack_1381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_321_delayed_4_0_337_inst_ack_1, ack => inputPort_1_Daemon_CP_1105_elements(91)); -- 
    -- CP-element group 92:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	60 
    -- CP-element group 92: 	91 
    -- CP-element group 92: 	72 
    -- CP-element group 92: marked-predecessors 
    -- CP-element group 92: 	94 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_3_341_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_3_341_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_3_341_Sample/req
      -- 
    req_1389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(92), ack => WPIPE_noblock_obuf_1_3_341_inst_req_0); -- 
    inputPort_1_Daemon_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_1105_elements(60) & inputPort_1_Daemon_CP_1105_elements(91) & inputPort_1_Daemon_CP_1105_elements(72) & inputPort_1_Daemon_CP_1105_elements(94);
      gj_inputPort_1_Daemon_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93: marked-successors 
    -- CP-element group 93: 	58 
    -- CP-element group 93: 	89 
    -- CP-element group 93: 	70 
    -- CP-element group 93:  members (6) 
      -- CP-element group 93: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_3_341_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_3_341_update_start_
      -- CP-element group 93: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_3_341_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_3_341_Sample/ack
      -- CP-element group 93: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_3_341_Update/$entry
      -- CP-element group 93: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_3_341_Update/req
      -- 
    ack_1390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_3_341_inst_ack_0, ack => inputPort_1_Daemon_CP_1105_elements(93)); -- 
    req_1394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(93), ack => WPIPE_noblock_obuf_1_3_341_inst_req_1); -- 
    -- CP-element group 94:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	102 
    -- CP-element group 94: marked-successors 
    -- CP-element group 94: 	92 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_3_341_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_3_341_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_3_341_Update/ack
      -- 
    ack_1395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_3_341_inst_ack_1, ack => inputPort_1_Daemon_CP_1105_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: marked-predecessors 
    -- CP-element group 95: 	99 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_346_update_start_
      -- CP-element group 95: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_346_Update/$entry
      -- CP-element group 95: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_346_Update/req
      -- 
    req_1408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(95), ack => W_data_to_outport_325_delayed_4_0_344_inst_req_1); -- 
    inputPort_1_Daemon_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_1_Daemon_CP_1105_elements(99);
      gj_inputPort_1_Daemon_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	38 
    -- CP-element group 96: successors 
    -- CP-element group 96: marked-successors 
    -- CP-element group 96: 	34 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_346_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_346_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_346_Sample/ack
      -- 
    ack_1404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_325_delayed_4_0_344_inst_ack_0, ack => inputPort_1_Daemon_CP_1105_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_346_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_346_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/assign_stmt_346_Update/ack
      -- 
    ack_1409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_325_delayed_4_0_344_inst_ack_1, ack => inputPort_1_Daemon_CP_1105_elements(97)); -- 
    -- CP-element group 98:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	60 
    -- CP-element group 98: 	97 
    -- CP-element group 98: 	76 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	100 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_4_348_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_4_348_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_4_348_Sample/req
      -- 
    req_1417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(98), ack => WPIPE_noblock_obuf_1_4_348_inst_req_0); -- 
    inputPort_1_Daemon_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_1105_elements(60) & inputPort_1_Daemon_CP_1105_elements(97) & inputPort_1_Daemon_CP_1105_elements(76) & inputPort_1_Daemon_CP_1105_elements(100);
      gj_inputPort_1_Daemon_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: marked-successors 
    -- CP-element group 99: 	58 
    -- CP-element group 99: 	95 
    -- CP-element group 99: 	74 
    -- CP-element group 99:  members (6) 
      -- CP-element group 99: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_4_348_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_4_348_update_start_
      -- CP-element group 99: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_4_348_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_4_348_Sample/ack
      -- CP-element group 99: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_4_348_Update/$entry
      -- CP-element group 99: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_4_348_Update/req
      -- 
    ack_1418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_4_348_inst_ack_0, ack => inputPort_1_Daemon_CP_1105_elements(99)); -- 
    req_1422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_1105_elements(99), ack => WPIPE_noblock_obuf_1_4_348_inst_req_1); -- 
    -- CP-element group 100:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100: marked-successors 
    -- CP-element group 100: 	98 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_4_348_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_4_348_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/WPIPE_noblock_obuf_1_4_348_Update/ack
      -- 
    ack_1423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_4_348_inst_ack_1, ack => inputPort_1_Daemon_CP_1105_elements(100)); -- 
    -- CP-element group 101:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	9 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	10 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group inputPort_1_Daemon_CP_1105_elements(101) is a control-delay.
    cp_element_101_delay: control_delay_element  generic map(name => " 101_delay", delay_value => 1)  port map(req => inputPort_1_Daemon_CP_1105_elements(9), ack => inputPort_1_Daemon_CP_1105_elements(101), clk => clk, reset =>reset);
    -- CP-element group 102:  join  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	12 
    -- CP-element group 102: 	13 
    -- CP-element group 102: 	88 
    -- CP-element group 102: 	94 
    -- CP-element group 102: 	100 
    -- CP-element group 102: 	82 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	6 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_214/do_while_stmt_215/do_while_stmt_215_loop_body/$exit
      -- 
    inputPort_1_Daemon_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 39) := "inputPort_1_Daemon_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_1105_elements(12) & inputPort_1_Daemon_CP_1105_elements(13) & inputPort_1_Daemon_CP_1105_elements(88) & inputPort_1_Daemon_CP_1105_elements(94) & inputPort_1_Daemon_CP_1105_elements(100) & inputPort_1_Daemon_CP_1105_elements(82);
      gj_inputPort_1_Daemon_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	5 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_214/do_while_stmt_215/loop_exit/$exit
      -- CP-element group 103: 	 branch_block_stmt_214/do_while_stmt_215/loop_exit/ack
      -- 
    ack_1428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_215_branch_ack_0, ack => inputPort_1_Daemon_CP_1105_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	5 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_214/do_while_stmt_215/loop_taken/$exit
      -- CP-element group 104: 	 branch_block_stmt_214/do_while_stmt_215/loop_taken/ack
      -- 
    ack_1432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_215_branch_ack_1, ack => inputPort_1_Daemon_CP_1105_elements(104)); -- 
    -- CP-element group 105:  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	3 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	1 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_214/do_while_stmt_215/$exit
      -- 
    inputPort_1_Daemon_CP_1105_elements(105) <= inputPort_1_Daemon_CP_1105_elements(3);
    inputPort_1_Daemon_do_while_stmt_215_terminator_1433: loop_terminator -- 
      generic map (name => " inputPort_1_Daemon_do_while_stmt_215_terminator_1433", max_iterations_in_flight =>7) 
      port map(loop_body_exit => inputPort_1_Daemon_CP_1105_elements(6),loop_continue => inputPort_1_Daemon_CP_1105_elements(104),loop_terminate => inputPort_1_Daemon_CP_1105_elements(103),loop_back => inputPort_1_Daemon_CP_1105_elements(4),loop_exit => inputPort_1_Daemon_CP_1105_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_217_phi_seq_1179_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_1_Daemon_CP_1105_elements(21);
      inputPort_1_Daemon_CP_1105_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_1_Daemon_CP_1105_elements(28);
      inputPort_1_Daemon_CP_1105_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_1_Daemon_CP_1105_elements(29);
      inputPort_1_Daemon_CP_1105_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_1_Daemon_CP_1105_elements(23);
      inputPort_1_Daemon_CP_1105_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_1_Daemon_CP_1105_elements(30);
      inputPort_1_Daemon_CP_1105_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_1_Daemon_CP_1105_elements(32);
      inputPort_1_Daemon_CP_1105_elements(24) <= phi_mux_reqs(1);
      phi_stmt_217_phi_seq_1179 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_217_phi_seq_1179") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_1_Daemon_CP_1105_elements(18), 
          phi_sample_ack => inputPort_1_Daemon_CP_1105_elements(19), 
          phi_update_req => inputPort_1_Daemon_CP_1105_elements(14), 
          phi_update_ack => inputPort_1_Daemon_CP_1105_elements(20), 
          phi_mux_ack => inputPort_1_Daemon_CP_1105_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_224_phi_seq_1241_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_1_Daemon_CP_1105_elements(44);
      inputPort_1_Daemon_CP_1105_elements(49)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_1_Daemon_CP_1105_elements(51);
      inputPort_1_Daemon_CP_1105_elements(50)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_1_Daemon_CP_1105_elements(52);
      inputPort_1_Daemon_CP_1105_elements(45) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_1_Daemon_CP_1105_elements(46);
      inputPort_1_Daemon_CP_1105_elements(53)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_1_Daemon_CP_1105_elements(53);
      inputPort_1_Daemon_CP_1105_elements(54)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_1_Daemon_CP_1105_elements(55);
      inputPort_1_Daemon_CP_1105_elements(47) <= phi_mux_reqs(1);
      phi_stmt_224_phi_seq_1241 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_224_phi_seq_1241") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_1_Daemon_CP_1105_elements(11), 
          phi_sample_ack => inputPort_1_Daemon_CP_1105_elements(41), 
          phi_update_req => inputPort_1_Daemon_CP_1105_elements(42), 
          phi_update_ack => inputPort_1_Daemon_CP_1105_elements(43), 
          phi_mux_ack => inputPort_1_Daemon_CP_1105_elements(48), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1130_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= inputPort_1_Daemon_CP_1105_elements(7);
        preds(1)  <= inputPort_1_Daemon_CP_1105_elements(8);
        entry_tmerge_1130 : transition_merge -- 
          generic map(name => " entry_tmerge_1130")
          port map (preds => preds, symbol_out => inputPort_1_Daemon_CP_1105_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal EQ_u8_u1_286_286_delayed_4_0_287 : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_293_293_delayed_4_0_297 : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_300_300_delayed_4_0_307 : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_307_307_delayed_4_0_317 : std_logic_vector(0 downto 0);
    signal RPIPE_in_data_1_223_wire : std_logic_vector(31 downto 0);
    signal R_ONE_1_270_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_16_220_wire_constant : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_257_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_260_wire : std_logic_vector(15 downto 0);
    signal SUB_u8_u8_278_wire : std_logic_vector(7 downto 0);
    signal continue_282 : std_logic_vector(0 downto 0);
    signal count_down_217 : std_logic_vector(15 downto 0);
    signal data_to_outport_273 : std_logic_vector(32 downto 0);
    signal data_to_outport_313_delayed_4_0_325 : std_logic_vector(32 downto 0);
    signal data_to_outport_317_delayed_4_0_332 : std_logic_vector(32 downto 0);
    signal data_to_outport_321_delayed_4_0_339 : std_logic_vector(32 downto 0);
    signal data_to_outport_325_delayed_4_0_346 : std_logic_vector(32 downto 0);
    signal dest_id_239 : std_logic_vector(7 downto 0);
    signal input_word_221 : std_logic_vector(31 downto 0);
    signal konst_227_wire_constant : std_logic_vector(7 downto 0);
    signal konst_233_wire_constant : std_logic_vector(15 downto 0);
    signal konst_256_wire_constant : std_logic_vector(15 downto 0);
    signal konst_259_wire_constant : std_logic_vector(15 downto 0);
    signal konst_275_wire_constant : std_logic_vector(7 downto 0);
    signal konst_277_wire_constant : std_logic_vector(7 downto 0);
    signal konst_285_wire_constant : std_logic_vector(7 downto 0);
    signal konst_295_wire_constant : std_logic_vector(7 downto 0);
    signal konst_305_wire_constant : std_logic_vector(7 downto 0);
    signal konst_315_wire_constant : std_logic_vector(7 downto 0);
    signal konst_362_wire_constant : std_logic_vector(0 downto 0);
    signal last_dest_id_224 : std_logic_vector(7 downto 0);
    signal new_packet_235 : std_logic_vector(0 downto 0);
    signal next_count_down_262 : std_logic_vector(15 downto 0);
    signal next_count_down_262_219_buffered : std_logic_vector(15 downto 0);
    signal next_last_dest_id_268 : std_logic_vector(7 downto 0);
    signal next_last_dest_id_268_226_buffered : std_logic_vector(7 downto 0);
    signal pkt_length_243 : std_logic_vector(15 downto 0);
    signal send_to_1_292 : std_logic_vector(0 downto 0);
    signal send_to_2_302 : std_logic_vector(0 downto 0);
    signal send_to_3_312 : std_logic_vector(0 downto 0);
    signal send_to_4_322 : std_logic_vector(0 downto 0);
    signal seq_id_247 : std_logic_vector(7 downto 0);
    signal type_cast_280_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_ONE_1_270_wire_constant <= "1";
    R_ZERO_16_220_wire_constant <= "0000000000000000";
    konst_227_wire_constant <= "00000000";
    konst_233_wire_constant <= "0000000000000000";
    konst_256_wire_constant <= "0000000000000001";
    konst_259_wire_constant <= "0000000000000001";
    konst_275_wire_constant <= "00000000";
    konst_277_wire_constant <= "00000001";
    konst_285_wire_constant <= "00000001";
    konst_295_wire_constant <= "00000010";
    konst_305_wire_constant <= "00000011";
    konst_315_wire_constant <= "00000100";
    konst_362_wire_constant <= "1";
    type_cast_280_wire_constant <= "1";
    phi_stmt_217: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= next_count_down_262_219_buffered & R_ZERO_16_220_wire_constant;
      req <= phi_stmt_217_req_0 & phi_stmt_217_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_217",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_217_ack_0,
          idata => idata,
          odata => count_down_217,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_217
    phi_stmt_224: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= next_last_dest_id_268_226_buffered & konst_227_wire_constant;
      req <= phi_stmt_224_req_0 & phi_stmt_224_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_224",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_224_ack_0,
          idata => idata,
          odata => last_dest_id_224,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_224
    -- flow-through select operator MUX_261_inst
    next_count_down_262 <= SUB_u16_u16_257_wire when (new_packet_235(0) /=  '0') else SUB_u16_u16_260_wire;
    -- flow-through select operator MUX_267_inst
    next_last_dest_id_268 <= dest_id_239 when (new_packet_235(0) /=  '0') else last_dest_id_224;
    -- flow-through slice operator slice_238_inst
    dest_id_239 <= input_word_221(31 downto 24);
    -- flow-through slice operator slice_242_inst
    pkt_length_243 <= input_word_221(23 downto 8);
    -- flow-through slice operator slice_246_inst
    seq_id_247 <= input_word_221(7 downto 0);
    W_data_to_outport_313_delayed_4_0_323_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_data_to_outport_313_delayed_4_0_323_inst_req_0;
      W_data_to_outport_313_delayed_4_0_323_inst_ack_0<= wack(0);
      rreq(0) <= W_data_to_outport_313_delayed_4_0_323_inst_req_1;
      W_data_to_outport_313_delayed_4_0_323_inst_ack_1<= rack(0);
      W_data_to_outport_313_delayed_4_0_323_inst : InterlockBuffer generic map ( -- 
        name => "W_data_to_outport_313_delayed_4_0_323_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 33,
        out_data_width => 33,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => data_to_outport_273,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => data_to_outport_313_delayed_4_0_325,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_data_to_outport_317_delayed_4_0_330_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_data_to_outport_317_delayed_4_0_330_inst_req_0;
      W_data_to_outport_317_delayed_4_0_330_inst_ack_0<= wack(0);
      rreq(0) <= W_data_to_outport_317_delayed_4_0_330_inst_req_1;
      W_data_to_outport_317_delayed_4_0_330_inst_ack_1<= rack(0);
      W_data_to_outport_317_delayed_4_0_330_inst : InterlockBuffer generic map ( -- 
        name => "W_data_to_outport_317_delayed_4_0_330_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 33,
        out_data_width => 33,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => data_to_outport_273,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => data_to_outport_317_delayed_4_0_332,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_data_to_outport_321_delayed_4_0_337_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_data_to_outport_321_delayed_4_0_337_inst_req_0;
      W_data_to_outport_321_delayed_4_0_337_inst_ack_0<= wack(0);
      rreq(0) <= W_data_to_outport_321_delayed_4_0_337_inst_req_1;
      W_data_to_outport_321_delayed_4_0_337_inst_ack_1<= rack(0);
      W_data_to_outport_321_delayed_4_0_337_inst : InterlockBuffer generic map ( -- 
        name => "W_data_to_outport_321_delayed_4_0_337_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 33,
        out_data_width => 33,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => data_to_outport_273,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => data_to_outport_321_delayed_4_0_339,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_data_to_outport_325_delayed_4_0_344_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_data_to_outport_325_delayed_4_0_344_inst_req_0;
      W_data_to_outport_325_delayed_4_0_344_inst_ack_0<= wack(0);
      rreq(0) <= W_data_to_outport_325_delayed_4_0_344_inst_req_1;
      W_data_to_outport_325_delayed_4_0_344_inst_ack_1<= rack(0);
      W_data_to_outport_325_delayed_4_0_344_inst : InterlockBuffer generic map ( -- 
        name => "W_data_to_outport_325_delayed_4_0_344_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 33,
        out_data_width => 33,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => data_to_outport_273,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => data_to_outport_325_delayed_4_0_346,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_count_down_262_219_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_count_down_262_219_buf_req_0;
      next_count_down_262_219_buf_ack_0<= wack(0);
      rreq(0) <= next_count_down_262_219_buf_req_1;
      next_count_down_262_219_buf_ack_1<= rack(0);
      next_count_down_262_219_buf : InterlockBuffer generic map ( -- 
        name => "next_count_down_262_219_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_count_down_262,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_count_down_262_219_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_last_dest_id_268_226_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_last_dest_id_268_226_buf_req_0;
      next_last_dest_id_268_226_buf_ack_0<= wack(0);
      rreq(0) <= next_last_dest_id_268_226_buf_req_1;
      next_last_dest_id_268_226_buf_ack_1<= rack(0);
      next_last_dest_id_268_226_buf : InterlockBuffer generic map ( -- 
        name => "next_last_dest_id_268_226_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_last_dest_id_268,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_last_dest_id_268_226_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_221
    process(RPIPE_in_data_1_223_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := RPIPE_in_data_1_223_wire(31 downto 0);
      input_word_221 <= tmp_var; -- 
    end process;
    do_while_stmt_215_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_362_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_215_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_215_branch_req_0,
          ack0 => do_while_stmt_215_branch_ack_0,
          ack1 => do_while_stmt_215_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- flow through binary operator AND_u1_u1_291_inst
    send_to_1_292 <= (EQ_u8_u1_286_286_delayed_4_0_287 and continue_282);
    -- flow through binary operator AND_u1_u1_301_inst
    send_to_2_302 <= (EQ_u8_u1_293_293_delayed_4_0_297 and continue_282);
    -- flow through binary operator AND_u1_u1_311_inst
    send_to_3_312 <= (EQ_u8_u1_300_300_delayed_4_0_307 and continue_282);
    -- flow through binary operator AND_u1_u1_321_inst
    send_to_4_322 <= (EQ_u8_u1_307_307_delayed_4_0_317 and continue_282);
    -- flow through binary operator CONCAT_u1_u33_272_inst
    process(R_ONE_1_270_wire_constant, input_word_221) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ONE_1_270_wire_constant, input_word_221, tmp_var);
      data_to_outport_273 <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u16_u1_234_inst
    process(count_down_217) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(count_down_217, konst_233_wire_constant, tmp_var);
      new_packet_235 <= tmp_var; --
    end process;
    -- shared split operator group (6) : EQ_u8_u1_286_inst 
    ApIntEq_group_6: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 4);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= next_last_dest_id_268;
      EQ_u8_u1_286_286_delayed_4_0_287 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u8_u1_286_inst_req_0;
      EQ_u8_u1_286_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u8_u1_286_inst_req_1;
      EQ_u8_u1_286_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_6_gI: SplitGuardInterface generic map(name => "ApIntEq_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000001",
          constant_width => 8,
          buffering  => 4,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : EQ_u8_u1_296_inst 
    ApIntEq_group_7: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 4);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= next_last_dest_id_268;
      EQ_u8_u1_293_293_delayed_4_0_297 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u8_u1_296_inst_req_0;
      EQ_u8_u1_296_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u8_u1_296_inst_req_1;
      EQ_u8_u1_296_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_7_gI: SplitGuardInterface generic map(name => "ApIntEq_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000010",
          constant_width => 8,
          buffering  => 4,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : EQ_u8_u1_306_inst 
    ApIntEq_group_8: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 4);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= next_last_dest_id_268;
      EQ_u8_u1_300_300_delayed_4_0_307 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u8_u1_306_inst_req_0;
      EQ_u8_u1_306_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u8_u1_306_inst_req_1;
      EQ_u8_u1_306_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_8_gI: SplitGuardInterface generic map(name => "ApIntEq_group_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_8",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000011",
          constant_width => 8,
          buffering  => 4,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : EQ_u8_u1_316_inst 
    ApIntEq_group_9: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 4);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= next_last_dest_id_268;
      EQ_u8_u1_307_307_delayed_4_0_317 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u8_u1_316_inst_req_0;
      EQ_u8_u1_316_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u8_u1_316_inst_req_1;
      EQ_u8_u1_316_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_9_gI: SplitGuardInterface generic map(name => "ApIntEq_group_9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_9",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000100",
          constant_width => 8,
          buffering  => 4,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- flow through binary operator SUB_u16_u16_257_inst
    SUB_u16_u16_257_wire <= std_logic_vector(unsigned(pkt_length_243) - unsigned(konst_256_wire_constant));
    -- flow through binary operator SUB_u16_u16_260_inst
    SUB_u16_u16_260_wire <= std_logic_vector(unsigned(count_down_217) - unsigned(konst_259_wire_constant));
    -- flow through binary operator SUB_u8_u8_278_inst
    SUB_u8_u8_278_wire <= std_logic_vector(unsigned(next_last_dest_id_268) - unsigned(konst_277_wire_constant));
    -- shared inport operator group (0) : RPIPE_in_data_1_223_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_in_data_1_223_inst_req_0;
      RPIPE_in_data_1_223_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_in_data_1_223_inst_req_1;
      RPIPE_in_data_1_223_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_in_data_1_223_wire <= data_out(31 downto 0);
      in_data_1_read_0_gI: SplitGuardInterface generic map(name => "in_data_1_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      in_data_1_read_0: InputPortRevised -- 
        generic map ( name => "in_data_1_read_0", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => in_data_1_pipe_read_req(0),
          oack => in_data_1_pipe_read_ack(0),
          odata => in_data_1_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_noblock_obuf_1_1_327_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_1_1_327_inst_req_0;
      WPIPE_noblock_obuf_1_1_327_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_1_1_327_inst_req_1;
      WPIPE_noblock_obuf_1_1_327_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_1_292(0);
      data_in <= data_to_outport_313_delayed_4_0_325;
      noblock_obuf_1_1_write_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_1_write_0: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_1_1", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_1_1_pipe_write_req(0),
          oack => noblock_obuf_1_1_pipe_write_ack(0),
          odata => noblock_obuf_1_1_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_noblock_obuf_1_2_334_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_1_2_334_inst_req_0;
      WPIPE_noblock_obuf_1_2_334_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_1_2_334_inst_req_1;
      WPIPE_noblock_obuf_1_2_334_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_2_302(0);
      data_in <= data_to_outport_317_delayed_4_0_332;
      noblock_obuf_1_2_write_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_2_write_1: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_1_2", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_1_2_pipe_write_req(0),
          oack => noblock_obuf_1_2_pipe_write_ack(0),
          odata => noblock_obuf_1_2_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_noblock_obuf_1_3_341_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_1_3_341_inst_req_0;
      WPIPE_noblock_obuf_1_3_341_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_1_3_341_inst_req_1;
      WPIPE_noblock_obuf_1_3_341_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_3_312(0);
      data_in <= data_to_outport_321_delayed_4_0_339;
      noblock_obuf_1_3_write_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_3_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_3_write_2: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_1_3", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_1_3_pipe_write_req(0),
          oack => noblock_obuf_1_3_pipe_write_ack(0),
          odata => noblock_obuf_1_3_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_noblock_obuf_1_4_348_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_1_4_348_inst_req_0;
      WPIPE_noblock_obuf_1_4_348_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_1_4_348_inst_req_1;
      WPIPE_noblock_obuf_1_4_348_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_4_322(0);
      data_in <= data_to_outport_325_delayed_4_0_346;
      noblock_obuf_1_4_write_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_4_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_4_write_3: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_1_4", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_1_4_pipe_write_req(0),
          oack => noblock_obuf_1_4_pipe_write_ack(0),
          odata => noblock_obuf_1_4_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared call operator group (0) : call_updateCounter_expr_281_inst 
    updateCounter_call_group_0: Block -- 
      signal data_in: std_logic_vector(16 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_updateCounter_expr_281_inst_req_0;
      call_updateCounter_expr_281_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_updateCounter_expr_281_inst_req_1;
      call_updateCounter_expr_281_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      updateCounter_call_group_0_gI: SplitGuardInterface generic map(name => "updateCounter_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_275_wire_constant & SUB_u8_u8_278_wire & type_cast_280_wire_constant;
      continue_282 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 17,
        owidth => 17,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => updateCounter_call_reqs(0),
          ackR => updateCounter_call_acks(0),
          dataR => updateCounter_call_data(16 downto 0),
          tagR => updateCounter_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => updateCounter_return_acks(0), -- cross-over
          ackL => updateCounter_return_reqs(0), -- cross-over
          dataL => updateCounter_return_data(0 downto 0),
          tagL => updateCounter_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end inputPort_1_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity inputPort_2_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    in_data_2_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_2_pipe_read_data : in   std_logic_vector(31 downto 0);
    noblock_obuf_2_1_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_1_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_2_2_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_2_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_2_3_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_3_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_2_4_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_4_pipe_write_data : out  std_logic_vector(32 downto 0);
    updateCounter_call_reqs : out  std_logic_vector(0 downto 0);
    updateCounter_call_acks : in   std_logic_vector(0 downto 0);
    updateCounter_call_data : out  std_logic_vector(16 downto 0);
    updateCounter_call_tag  :  out  std_logic_vector(0 downto 0);
    updateCounter_return_reqs : out  std_logic_vector(0 downto 0);
    updateCounter_return_acks : in   std_logic_vector(0 downto 0);
    updateCounter_return_data : in   std_logic_vector(0 downto 0);
    updateCounter_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity inputPort_2_Daemon;
architecture inputPort_2_Daemon_arch of inputPort_2_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal inputPort_2_Daemon_CP_1434_start: Boolean;
  signal inputPort_2_Daemon_CP_1434_symbol: Boolean;
  -- volatile/operator module components. 
  component updateCounter is -- 
    generic (tag_length : integer); 
    port ( -- 
      input_port : in  std_logic_vector(7 downto 0);
      output_port : in  std_logic_vector(7 downto 0);
      up : in  std_logic_vector(0 downto 0);
      continue : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(3 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(1 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(1 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal EQ_u8_u1_438_inst_ack_1 : boolean;
  signal EQ_u8_u1_448_inst_req_1 : boolean;
  signal EQ_u8_u1_438_inst_ack_0 : boolean;
  signal EQ_u8_u1_458_inst_ack_0 : boolean;
  signal RPIPE_in_data_2_375_inst_req_1 : boolean;
  signal EQ_u8_u1_438_inst_req_1 : boolean;
  signal do_while_stmt_367_branch_req_0 : boolean;
  signal next_last_dest_id_420_379_buf_req_0 : boolean;
  signal call_updateCounter_expr_433_inst_req_0 : boolean;
  signal phi_stmt_369_req_1 : boolean;
  signal next_count_down_414_372_buf_req_1 : boolean;
  signal phi_stmt_369_req_0 : boolean;
  signal RPIPE_in_data_2_375_inst_ack_1 : boolean;
  signal next_count_down_414_372_buf_ack_0 : boolean;
  signal next_count_down_414_372_buf_req_0 : boolean;
  signal EQ_u8_u1_448_inst_ack_1 : boolean;
  signal call_updateCounter_expr_433_inst_ack_1 : boolean;
  signal phi_stmt_369_ack_0 : boolean;
  signal W_data_to_outport_445_delayed_4_0_482_inst_req_0 : boolean;
  signal EQ_u8_u1_458_inst_req_1 : boolean;
  signal EQ_u8_u1_448_inst_ack_0 : boolean;
  signal W_data_to_outport_441_delayed_4_0_475_inst_ack_1 : boolean;
  signal EQ_u8_u1_458_inst_ack_1 : boolean;
  signal phi_stmt_376_req_1 : boolean;
  signal WPIPE_noblock_obuf_2_1_479_inst_ack_1 : boolean;
  signal EQ_u8_u1_468_inst_ack_1 : boolean;
  signal call_updateCounter_expr_433_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_2_3_493_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_2_3_493_inst_ack_1 : boolean;
  signal next_count_down_414_372_buf_ack_1 : boolean;
  signal W_data_to_outport_449_delayed_4_0_489_inst_req_0 : boolean;
  signal W_data_to_outport_449_delayed_4_0_489_inst_ack_0 : boolean;
  signal W_data_to_outport_453_delayed_4_0_496_inst_ack_1 : boolean;
  signal EQ_u8_u1_458_inst_req_0 : boolean;
  signal W_data_to_outport_449_delayed_4_0_489_inst_req_1 : boolean;
  signal W_data_to_outport_449_delayed_4_0_489_inst_ack_1 : boolean;
  signal call_updateCounter_expr_433_inst_req_1 : boolean;
  signal next_last_dest_id_420_379_buf_ack_0 : boolean;
  signal WPIPE_noblock_obuf_2_3_493_inst_ack_0 : boolean;
  signal EQ_u8_u1_468_inst_req_0 : boolean;
  signal EQ_u8_u1_468_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_2_4_500_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_2_4_500_inst_req_1 : boolean;
  signal do_while_stmt_367_branch_ack_0 : boolean;
  signal WPIPE_noblock_obuf_2_4_500_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_2_4_500_inst_ack_0 : boolean;
  signal phi_stmt_376_req_0 : boolean;
  signal RPIPE_in_data_2_375_inst_ack_0 : boolean;
  signal EQ_u8_u1_438_inst_req_0 : boolean;
  signal EQ_u8_u1_448_inst_req_0 : boolean;
  signal EQ_u8_u1_468_inst_req_1 : boolean;
  signal RPIPE_in_data_2_375_inst_req_0 : boolean;
  signal next_last_dest_id_420_379_buf_ack_1 : boolean;
  signal phi_stmt_376_ack_0 : boolean;
  signal next_last_dest_id_420_379_buf_req_1 : boolean;
  signal W_data_to_outport_441_delayed_4_0_475_inst_req_1 : boolean;
  signal W_data_to_outport_445_delayed_4_0_482_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_2_2_486_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_2_2_486_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_2_2_486_inst_req_0 : boolean;
  signal W_data_to_outport_441_delayed_4_0_475_inst_ack_0 : boolean;
  signal W_data_to_outport_441_delayed_4_0_475_inst_req_0 : boolean;
  signal W_data_to_outport_445_delayed_4_0_482_inst_ack_1 : boolean;
  signal W_data_to_outport_445_delayed_4_0_482_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_2_1_479_inst_ack_0 : boolean;
  signal W_data_to_outport_453_delayed_4_0_496_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_2_2_486_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_2_3_493_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_2_1_479_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_2_1_479_inst_req_1 : boolean;
  signal W_data_to_outport_453_delayed_4_0_496_inst_req_0 : boolean;
  signal W_data_to_outport_453_delayed_4_0_496_inst_ack_0 : boolean;
  signal do_while_stmt_367_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "inputPort_2_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  inputPort_2_Daemon_CP_1434_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "inputPort_2_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_2_Daemon_CP_1434_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= inputPort_2_Daemon_CP_1434_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_2_Daemon_CP_1434_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  inputPort_2_Daemon_CP_1434: Block -- control-path 
    signal inputPort_2_Daemon_CP_1434_elements: BooleanArray(105 downto 0);
    -- 
  begin -- 
    inputPort_2_Daemon_CP_1434_elements(0) <= inputPort_2_Daemon_CP_1434_start;
    inputPort_2_Daemon_CP_1434_symbol <= inputPort_2_Daemon_CP_1434_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_366/do_while_stmt_367__entry__
      -- CP-element group 0: 	 branch_block_stmt_366/branch_block_stmt_366__entry__
      -- CP-element group 0: 	 branch_block_stmt_366/$entry
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	105 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_366/do_while_stmt_367__exit__
      -- CP-element group 1: 	 branch_block_stmt_366/branch_block_stmt_366__exit__
      -- CP-element group 1: 	 branch_block_stmt_366/$exit
      -- CP-element group 1: 	 $exit
      -- 
    inputPort_2_Daemon_CP_1434_elements(1) <= inputPort_2_Daemon_CP_1434_elements(105);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367__entry__
      -- CP-element group 2: 	 branch_block_stmt_366/do_while_stmt_367/$entry
      -- 
    inputPort_2_Daemon_CP_1434_elements(2) <= inputPort_2_Daemon_CP_1434_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	105 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367__exit__
      -- 
    -- Element group inputPort_2_Daemon_CP_1434_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_366/do_while_stmt_367/loop_back
      -- 
    -- Element group inputPort_2_Daemon_CP_1434_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	103 
    -- CP-element group 5: 	104 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_366/do_while_stmt_367/condition_done
      -- CP-element group 5: 	 branch_block_stmt_366/do_while_stmt_367/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_366/do_while_stmt_367/loop_taken/$entry
      -- 
    inputPort_2_Daemon_CP_1434_elements(5) <= inputPort_2_Daemon_CP_1434_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	102 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_366/do_while_stmt_367/loop_body_done
      -- 
    inputPort_2_Daemon_CP_1434_elements(6) <= inputPort_2_Daemon_CP_1434_elements(102);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	20 
    -- CP-element group 7: 	44 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/back_edge_to_loop_body
      -- 
    inputPort_2_Daemon_CP_1434_elements(7) <= inputPort_2_Daemon_CP_1434_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	22 
    -- CP-element group 8: 	46 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/first_time_through_loop_body
      -- 
    inputPort_2_Daemon_CP_1434_elements(8) <= inputPort_2_Daemon_CP_1434_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	17 
    -- CP-element group 9: 	101 
    -- CP-element group 9: 	33 
    -- CP-element group 9: 	38 
    -- CP-element group 9: 	39 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_373_sample_start_
      -- 
    -- Element group inputPort_2_Daemon_CP_1434_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	101 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/condition_evaluated
      -- 
    condition_evaluated_1458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(10), ack => do_while_stmt_367_branch_req_0); -- 
    inputPort_2_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_1434_elements(15) & inputPort_2_Daemon_CP_1434_elements(101);
      gj_inputPort_2_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	16 
    -- CP-element group 11: 	38 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	40 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_369_sample_start__ps
      -- 
    inputPort_2_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_1434_elements(9) & inputPort_2_Daemon_CP_1434_elements(16) & inputPort_2_Daemon_CP_1434_elements(38) & inputPort_2_Daemon_CP_1434_elements(15);
      gj_inputPort_2_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	18 
    -- CP-element group 12: 	36 
    -- CP-element group 12: 	41 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12: 	102 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	16 
    -- CP-element group 12: 	38 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_369_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_376_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_373_sample_completed_
      -- 
    inputPort_2_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_1434_elements(18) & inputPort_2_Daemon_CP_1434_elements(36) & inputPort_2_Daemon_CP_1434_elements(41);
      gj_inputPort_2_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	102 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/aggregated_phi_sample_ack_d
      -- 
    -- Element group inputPort_2_Daemon_CP_1434_elements(13) is a control-delay.
    cp_element_13_delay: control_delay_element  generic map(name => " 13_delay", delay_value => 1)  port map(req => inputPort_2_Daemon_CP_1434_elements(12), ack => inputPort_2_Daemon_CP_1434_elements(13), clk => clk, reset =>reset);
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	17 
    -- CP-element group 14: 	33 
    -- CP-element group 14: 	39 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	35 
    -- CP-element group 14: 	42 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/aggregated_phi_update_req
      -- CP-element group 14: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_369_update_start__ps
      -- 
    inputPort_2_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_1434_elements(17) & inputPort_2_Daemon_CP_1434_elements(33) & inputPort_2_Daemon_CP_1434_elements(39);
      gj_inputPort_2_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	19 
    -- CP-element group 15: 	37 
    -- CP-element group 15: 	43 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/aggregated_phi_update_ack
      -- 
    inputPort_2_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_1434_elements(19) & inputPort_2_Daemon_CP_1434_elements(37) & inputPort_2_Daemon_CP_1434_elements(43);
      gj_inputPort_2_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	11 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_369_sample_start_
      -- 
    inputPort_2_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_1434_elements(9) & inputPort_2_Daemon_CP_1434_elements(12);
      gj_inputPort_2_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	9 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	67 
    -- CP-element group 17: 	71 
    -- CP-element group 17: 	75 
    -- CP-element group 17: 	63 
    -- CP-element group 17: 	59 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	14 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_369_update_start_
      -- 
    inputPort_2_Daemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_1434_elements(9) & inputPort_2_Daemon_CP_1434_elements(67) & inputPort_2_Daemon_CP_1434_elements(71) & inputPort_2_Daemon_CP_1434_elements(75) & inputPort_2_Daemon_CP_1434_elements(63) & inputPort_2_Daemon_CP_1434_elements(59);
      gj_inputPort_2_Daemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_369_sample_completed__ps
      -- 
    -- Element group inputPort_2_Daemon_CP_1434_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: 	65 
    -- CP-element group 19: 	69 
    -- CP-element group 19: 	73 
    -- CP-element group 19: 	61 
    -- CP-element group 19: 	57 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_369_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_369_update_completed__ps
      -- 
    -- Element group inputPort_2_Daemon_CP_1434_elements(19) is bound as output of CP function.
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	7 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_369_loopback_trigger
      -- 
    inputPort_2_Daemon_CP_1434_elements(20) <= inputPort_2_Daemon_CP_1434_elements(7);
    -- CP-element group 21:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_369_loopback_sample_req
      -- CP-element group 21: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_369_loopback_sample_req_ps
      -- 
    phi_stmt_369_loopback_sample_req_1474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_369_loopback_sample_req_1474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(21), ack => phi_stmt_369_req_1); -- 
    -- Element group inputPort_2_Daemon_CP_1434_elements(21) is bound as output of CP function.
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	8 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_369_entry_trigger
      -- 
    inputPort_2_Daemon_CP_1434_elements(22) <= inputPort_2_Daemon_CP_1434_elements(8);
    -- CP-element group 23:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_369_entry_sample_req_ps
      -- CP-element group 23: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_369_entry_sample_req
      -- 
    phi_stmt_369_entry_sample_req_1477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_369_entry_sample_req_1477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(23), ack => phi_stmt_369_req_0); -- 
    -- Element group inputPort_2_Daemon_CP_1434_elements(23) is bound as output of CP function.
    -- CP-element group 24:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_369_phi_mux_ack
      -- CP-element group 24: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_369_phi_mux_ack_ps
      -- 
    phi_stmt_369_phi_mux_ack_1480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_369_ack_0, ack => inputPort_2_Daemon_CP_1434_elements(24)); -- 
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_ZERO_16_371_sample_start__ps
      -- CP-element group 25: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_ZERO_16_371_sample_completed__ps
      -- CP-element group 25: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_ZERO_16_371_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_ZERO_16_371_sample_start_
      -- 
    -- Element group inputPort_2_Daemon_CP_1434_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_ZERO_16_371_update_start__ps
      -- CP-element group 26: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_ZERO_16_371_update_start_
      -- 
    -- Element group inputPort_2_Daemon_CP_1434_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	28 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_ZERO_16_371_update_completed__ps
      -- 
    inputPort_2_Daemon_CP_1434_elements(27) <= inputPort_2_Daemon_CP_1434_elements(28);
    -- CP-element group 28:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	27 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_ZERO_16_371_update_completed_
      -- 
    -- Element group inputPort_2_Daemon_CP_1434_elements(28) is a control-delay.
    cp_element_28_delay: control_delay_element  generic map(name => " 28_delay", delay_value => 1)  port map(req => inputPort_2_Daemon_CP_1434_elements(26), ack => inputPort_2_Daemon_CP_1434_elements(28), clk => clk, reset =>reset);
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_count_down_372_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_count_down_372_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_count_down_372_Sample/req
      -- CP-element group 29: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_count_down_372_sample_start__ps
      -- 
    req_1501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(29), ack => next_count_down_414_372_buf_req_0); -- 
    -- Element group inputPort_2_Daemon_CP_1434_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_count_down_372_Update/req
      -- CP-element group 30: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_count_down_372_update_start__ps
      -- CP-element group 30: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_count_down_372_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_count_down_372_update_start_
      -- 
    req_1506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(30), ack => next_count_down_414_372_buf_req_1); -- 
    -- Element group inputPort_2_Daemon_CP_1434_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_count_down_372_Sample/ack
      -- CP-element group 31: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_count_down_372_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_count_down_372_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_count_down_372_sample_completed__ps
      -- 
    ack_1502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_414_372_buf_ack_0, ack => inputPort_2_Daemon_CP_1434_elements(31)); -- 
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_count_down_372_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_count_down_372_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_count_down_372_update_completed__ps
      -- CP-element group 32: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_count_down_372_Update/ack
      -- 
    ack_1507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_414_372_buf_ack_1, ack => inputPort_2_Daemon_CP_1434_elements(32)); -- 
    -- CP-element group 33:  join  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	9 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	84 
    -- CP-element group 33: 	90 
    -- CP-element group 33: 	96 
    -- CP-element group 33: 	67 
    -- CP-element group 33: 	71 
    -- CP-element group 33: 	75 
    -- CP-element group 33: 	63 
    -- CP-element group 33: 	78 
    -- CP-element group 33: 	59 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	14 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_373_update_start_
      -- 
    inputPort_2_Daemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_1434_elements(9) & inputPort_2_Daemon_CP_1434_elements(84) & inputPort_2_Daemon_CP_1434_elements(90) & inputPort_2_Daemon_CP_1434_elements(96) & inputPort_2_Daemon_CP_1434_elements(67) & inputPort_2_Daemon_CP_1434_elements(71) & inputPort_2_Daemon_CP_1434_elements(75) & inputPort_2_Daemon_CP_1434_elements(63) & inputPort_2_Daemon_CP_1434_elements(78) & inputPort_2_Daemon_CP_1434_elements(59);
      gj_inputPort_2_Daemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	11 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	37 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/RPIPE_in_data_2_375_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/RPIPE_in_data_2_375_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/RPIPE_in_data_2_375_Sample/$entry
      -- 
    rr_1520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(34), ack => RPIPE_in_data_2_375_inst_req_0); -- 
    inputPort_2_Daemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_1434_elements(11) & inputPort_2_Daemon_CP_1434_elements(37);
      gj_inputPort_2_Daemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	14 
    -- CP-element group 35: 	36 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/RPIPE_in_data_2_375_Update/cr
      -- CP-element group 35: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/RPIPE_in_data_2_375_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/RPIPE_in_data_2_375_update_start_
      -- 
    cr_1525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(35), ack => RPIPE_in_data_2_375_inst_req_1); -- 
    inputPort_2_Daemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_1434_elements(14) & inputPort_2_Daemon_CP_1434_elements(36);
      gj_inputPort_2_Daemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	12 
    -- CP-element group 36: 	35 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/RPIPE_in_data_2_375_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/RPIPE_in_data_2_375_Sample/ra
      -- CP-element group 36: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/RPIPE_in_data_2_375_Sample/$exit
      -- 
    ra_1521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_2_375_inst_ack_0, ack => inputPort_2_Daemon_CP_1434_elements(36)); -- 
    -- CP-element group 37:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	84 
    -- CP-element group 37: 	15 
    -- CP-element group 37: 	90 
    -- CP-element group 37: 	96 
    -- CP-element group 37: 	65 
    -- CP-element group 37: 	69 
    -- CP-element group 37: 	73 
    -- CP-element group 37: 	61 
    -- CP-element group 37: 	78 
    -- CP-element group 37: 	57 
    -- CP-element group 37: marked-successors 
    -- CP-element group 37: 	34 
    -- CP-element group 37:  members (16) 
      -- CP-element group 37: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/RPIPE_in_data_2_375_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_373_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/RPIPE_in_data_2_375_Update/ca
      -- CP-element group 37: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/RPIPE_in_data_2_375_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_484_Sample/req
      -- CP-element group 37: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_491_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_491_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_491_Sample/req
      -- CP-element group 37: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_477_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_477_Sample/req
      -- CP-element group 37: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_477_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_484_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_498_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_484_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_498_Sample/req
      -- CP-element group 37: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_498_sample_start_
      -- 
    ca_1526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_2_375_inst_ack_1, ack => inputPort_2_Daemon_CP_1434_elements(37)); -- 
    req_1676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(37), ack => W_data_to_outport_445_delayed_4_0_482_inst_req_0); -- 
    req_1704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(37), ack => W_data_to_outport_449_delayed_4_0_489_inst_req_0); -- 
    req_1732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(37), ack => W_data_to_outport_453_delayed_4_0_496_inst_req_0); -- 
    req_1648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(37), ack => W_data_to_outport_441_delayed_4_0_475_inst_req_0); -- 
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	9 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	12 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	11 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_376_sample_start_
      -- 
    inputPort_2_Daemon_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_1434_elements(9) & inputPort_2_Daemon_CP_1434_elements(12);
      gj_inputPort_2_Daemon_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  join  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	9 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	67 
    -- CP-element group 39: 	71 
    -- CP-element group 39: 	75 
    -- CP-element group 39: 	63 
    -- CP-element group 39: 	59 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	14 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_376_update_start_
      -- 
    inputPort_2_Daemon_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_1434_elements(9) & inputPort_2_Daemon_CP_1434_elements(67) & inputPort_2_Daemon_CP_1434_elements(71) & inputPort_2_Daemon_CP_1434_elements(75) & inputPort_2_Daemon_CP_1434_elements(63) & inputPort_2_Daemon_CP_1434_elements(59);
      gj_inputPort_2_Daemon_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	11 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_376_sample_start__ps
      -- 
    inputPort_2_Daemon_CP_1434_elements(40) <= inputPort_2_Daemon_CP_1434_elements(11);
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	12 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_376_sample_completed__ps
      -- 
    -- Element group inputPort_2_Daemon_CP_1434_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	14 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_376_update_start__ps
      -- 
    inputPort_2_Daemon_CP_1434_elements(42) <= inputPort_2_Daemon_CP_1434_elements(14);
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	15 
    -- CP-element group 43: 	65 
    -- CP-element group 43: 	69 
    -- CP-element group 43: 	73 
    -- CP-element group 43: 	61 
    -- CP-element group 43: 	57 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_376_update_completed__ps
      -- CP-element group 43: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_376_update_completed_
      -- 
    -- Element group inputPort_2_Daemon_CP_1434_elements(43) is bound as output of CP function.
    -- CP-element group 44:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	7 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_376_loopback_trigger
      -- 
    inputPort_2_Daemon_CP_1434_elements(44) <= inputPort_2_Daemon_CP_1434_elements(7);
    -- CP-element group 45:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_376_loopback_sample_req
      -- CP-element group 45: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_376_loopback_sample_req_ps
      -- 
    phi_stmt_376_loopback_sample_req_1536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_376_loopback_sample_req_1536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(45), ack => phi_stmt_376_req_1); -- 
    -- Element group inputPort_2_Daemon_CP_1434_elements(45) is bound as output of CP function.
    -- CP-element group 46:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	8 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_376_entry_trigger
      -- 
    inputPort_2_Daemon_CP_1434_elements(46) <= inputPort_2_Daemon_CP_1434_elements(8);
    -- CP-element group 47:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_376_entry_sample_req_ps
      -- CP-element group 47: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_376_entry_sample_req
      -- 
    phi_stmt_376_entry_sample_req_1539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_376_entry_sample_req_1539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(47), ack => phi_stmt_376_req_0); -- 
    -- Element group inputPort_2_Daemon_CP_1434_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_376_phi_mux_ack_ps
      -- CP-element group 48: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/phi_stmt_376_phi_mux_ack
      -- 
    phi_stmt_376_phi_mux_ack_1542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_376_ack_0, ack => inputPort_2_Daemon_CP_1434_elements(48)); -- 
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/konst_378_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/konst_378_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/konst_378_sample_completed__ps
      -- CP-element group 49: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/konst_378_sample_start__ps
      -- 
    -- Element group inputPort_2_Daemon_CP_1434_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (2) 
      -- CP-element group 50: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/konst_378_update_start_
      -- CP-element group 50: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/konst_378_update_start__ps
      -- 
    -- Element group inputPort_2_Daemon_CP_1434_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	52 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/konst_378_update_completed__ps
      -- 
    inputPort_2_Daemon_CP_1434_elements(51) <= inputPort_2_Daemon_CP_1434_elements(52);
    -- CP-element group 52:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	51 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/konst_378_update_completed_
      -- 
    -- Element group inputPort_2_Daemon_CP_1434_elements(52) is a control-delay.
    cp_element_52_delay: control_delay_element  generic map(name => " 52_delay", delay_value => 1)  port map(req => inputPort_2_Daemon_CP_1434_elements(50), ack => inputPort_2_Daemon_CP_1434_elements(52), clk => clk, reset =>reset);
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_last_dest_id_379_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_last_dest_id_379_Sample/req
      -- CP-element group 53: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_last_dest_id_379_sample_start__ps
      -- CP-element group 53: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_last_dest_id_379_sample_start_
      -- 
    req_1563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(53), ack => next_last_dest_id_420_379_buf_req_0); -- 
    -- Element group inputPort_2_Daemon_CP_1434_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_last_dest_id_379_update_start_
      -- CP-element group 54: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_last_dest_id_379_Update/req
      -- CP-element group 54: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_last_dest_id_379_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_last_dest_id_379_update_start__ps
      -- 
    req_1568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(54), ack => next_last_dest_id_420_379_buf_req_1); -- 
    -- Element group inputPort_2_Daemon_CP_1434_elements(54) is bound as output of CP function.
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_last_dest_id_379_sample_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_last_dest_id_379_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_last_dest_id_379_Sample/ack
      -- CP-element group 55: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_last_dest_id_379_sample_completed_
      -- 
    ack_1564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_420_379_buf_ack_0, ack => inputPort_2_Daemon_CP_1434_elements(55)); -- 
    -- CP-element group 56:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_last_dest_id_379_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_last_dest_id_379_Update/ack
      -- CP-element group 56: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_last_dest_id_379_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/R_next_last_dest_id_379_update_completed__ps
      -- 
    ack_1569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_420_379_buf_ack_1, ack => inputPort_2_Daemon_CP_1434_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	19 
    -- CP-element group 57: 	37 
    -- CP-element group 57: 	43 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/call_updateCounter_expr_433_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/call_updateCounter_expr_433_Sample/req
      -- CP-element group 57: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/call_updateCounter_expr_433_sample_start_
      -- 
    req_1578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(57), ack => call_updateCounter_expr_433_inst_req_0); -- 
    inputPort_2_Daemon_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_1434_elements(19) & inputPort_2_Daemon_CP_1434_elements(37) & inputPort_2_Daemon_CP_1434_elements(43);
      gj_inputPort_2_Daemon_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	81 
    -- CP-element group 58: 	87 
    -- CP-element group 58: 	93 
    -- CP-element group 58: 	99 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/call_updateCounter_expr_433_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/call_updateCounter_expr_433_Update/req
      -- CP-element group 58: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/call_updateCounter_expr_433_update_start_
      -- 
    req_1583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(58), ack => call_updateCounter_expr_433_inst_req_1); -- 
    inputPort_2_Daemon_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_1434_elements(81) & inputPort_2_Daemon_CP_1434_elements(87) & inputPort_2_Daemon_CP_1434_elements(93) & inputPort_2_Daemon_CP_1434_elements(99);
      gj_inputPort_2_Daemon_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: marked-successors 
    -- CP-element group 59: 	17 
    -- CP-element group 59: 	33 
    -- CP-element group 59: 	39 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/call_updateCounter_expr_433_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/call_updateCounter_expr_433_Sample/ack
      -- CP-element group 59: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/call_updateCounter_expr_433_sample_completed_
      -- 
    ack_1579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_updateCounter_expr_433_inst_ack_0, ack => inputPort_2_Daemon_CP_1434_elements(59)); -- 
    -- CP-element group 60:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	80 
    -- CP-element group 60: 	86 
    -- CP-element group 60: 	92 
    -- CP-element group 60: 	98 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/call_updateCounter_expr_433_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/call_updateCounter_expr_433_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/call_updateCounter_expr_433_update_completed_
      -- 
    ack_1584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_updateCounter_expr_433_inst_ack_1, ack => inputPort_2_Daemon_CP_1434_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	19 
    -- CP-element group 61: 	37 
    -- CP-element group 61: 	43 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_438_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_438_Sample/rr
      -- CP-element group 61: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_438_Sample/$entry
      -- 
    rr_1592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(61), ack => EQ_u8_u1_438_inst_req_0); -- 
    inputPort_2_Daemon_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_1434_elements(19) & inputPort_2_Daemon_CP_1434_elements(37) & inputPort_2_Daemon_CP_1434_elements(43);
      gj_inputPort_2_Daemon_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	81 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_438_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_438_Update/cr
      -- CP-element group 62: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_438_update_start_
      -- 
    cr_1597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(62), ack => EQ_u8_u1_438_inst_req_1); -- 
    inputPort_2_Daemon_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_2_Daemon_CP_1434_elements(81);
      gj_inputPort_2_Daemon_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	17 
    -- CP-element group 63: 	33 
    -- CP-element group 63: 	39 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_438_Sample/ra
      -- CP-element group 63: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_438_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_438_Sample/$exit
      -- 
    ra_1593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_438_inst_ack_0, ack => inputPort_2_Daemon_CP_1434_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	80 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_438_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_438_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_438_update_completed_
      -- 
    ca_1598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_438_inst_ack_1, ack => inputPort_2_Daemon_CP_1434_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	19 
    -- CP-element group 65: 	37 
    -- CP-element group 65: 	43 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_448_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_448_Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_448_Sample/$entry
      -- 
    rr_1606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(65), ack => EQ_u8_u1_448_inst_req_0); -- 
    inputPort_2_Daemon_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_1434_elements(19) & inputPort_2_Daemon_CP_1434_elements(37) & inputPort_2_Daemon_CP_1434_elements(43);
      gj_inputPort_2_Daemon_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	87 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_448_Update/cr
      -- CP-element group 66: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_448_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_448_update_start_
      -- 
    cr_1611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(66), ack => EQ_u8_u1_448_inst_req_1); -- 
    inputPort_2_Daemon_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_2_Daemon_CP_1434_elements(87);
      gj_inputPort_2_Daemon_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	17 
    -- CP-element group 67: 	33 
    -- CP-element group 67: 	39 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_448_Sample/ra
      -- CP-element group 67: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_448_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_448_Sample/$exit
      -- 
    ra_1607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_448_inst_ack_0, ack => inputPort_2_Daemon_CP_1434_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	86 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_448_Update/ca
      -- CP-element group 68: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_448_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_448_update_completed_
      -- 
    ca_1612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_448_inst_ack_1, ack => inputPort_2_Daemon_CP_1434_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	19 
    -- CP-element group 69: 	37 
    -- CP-element group 69: 	43 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_458_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_458_Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_458_sample_start_
      -- 
    rr_1620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(69), ack => EQ_u8_u1_458_inst_req_0); -- 
    inputPort_2_Daemon_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_1434_elements(19) & inputPort_2_Daemon_CP_1434_elements(37) & inputPort_2_Daemon_CP_1434_elements(43);
      gj_inputPort_2_Daemon_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	93 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_458_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_458_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_458_update_start_
      -- 
    cr_1625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(70), ack => EQ_u8_u1_458_inst_req_1); -- 
    inputPort_2_Daemon_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_2_Daemon_CP_1434_elements(93);
      gj_inputPort_2_Daemon_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: marked-successors 
    -- CP-element group 71: 	17 
    -- CP-element group 71: 	33 
    -- CP-element group 71: 	39 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_458_Sample/ra
      -- CP-element group 71: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_458_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_458_sample_completed_
      -- 
    ra_1621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_458_inst_ack_0, ack => inputPort_2_Daemon_CP_1434_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	92 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_458_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_458_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_458_update_completed_
      -- 
    ca_1626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_458_inst_ack_1, ack => inputPort_2_Daemon_CP_1434_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	19 
    -- CP-element group 73: 	37 
    -- CP-element group 73: 	43 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_468_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_468_Sample/rr
      -- CP-element group 73: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_468_Sample/$entry
      -- 
    rr_1634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(73), ack => EQ_u8_u1_468_inst_req_0); -- 
    inputPort_2_Daemon_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_1434_elements(19) & inputPort_2_Daemon_CP_1434_elements(37) & inputPort_2_Daemon_CP_1434_elements(43);
      gj_inputPort_2_Daemon_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	99 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_468_update_start_
      -- CP-element group 74: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_468_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_468_Update/cr
      -- 
    cr_1639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(74), ack => EQ_u8_u1_468_inst_req_1); -- 
    inputPort_2_Daemon_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_2_Daemon_CP_1434_elements(99);
      gj_inputPort_2_Daemon_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	17 
    -- CP-element group 75: 	33 
    -- CP-element group 75: 	39 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_468_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_468_Sample/ra
      -- CP-element group 75: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_468_Sample/$exit
      -- 
    ra_1635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_468_inst_ack_0, ack => inputPort_2_Daemon_CP_1434_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	98 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_468_Update/ca
      -- CP-element group 76: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_468_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/EQ_u8_u1_468_Update/$exit
      -- 
    ca_1640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_468_inst_ack_1, ack => inputPort_2_Daemon_CP_1434_elements(76)); -- 
    -- CP-element group 77:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	81 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_477_update_start_
      -- CP-element group 77: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_477_Update/req
      -- CP-element group 77: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_477_Update/$entry
      -- 
    req_1653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(77), ack => W_data_to_outport_441_delayed_4_0_475_inst_req_1); -- 
    inputPort_2_Daemon_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_2_Daemon_CP_1434_elements(81);
      gj_inputPort_2_Daemon_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	37 
    -- CP-element group 78: successors 
    -- CP-element group 78: marked-successors 
    -- CP-element group 78: 	33 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_477_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_477_Sample/ack
      -- CP-element group 78: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_477_Sample/$exit
      -- 
    ack_1649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_441_delayed_4_0_475_inst_ack_0, ack => inputPort_2_Daemon_CP_1434_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_477_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_477_Update/ack
      -- CP-element group 79: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_477_update_completed_
      -- 
    ack_1654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_441_delayed_4_0_475_inst_ack_1, ack => inputPort_2_Daemon_CP_1434_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: 	60 
    -- CP-element group 80: 	64 
    -- CP-element group 80: marked-predecessors 
    -- CP-element group 80: 	82 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_1_479_Sample/req
      -- CP-element group 80: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_1_479_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_1_479_sample_start_
      -- 
    req_1662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(80), ack => WPIPE_noblock_obuf_2_1_479_inst_req_0); -- 
    inputPort_2_Daemon_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_1434_elements(79) & inputPort_2_Daemon_CP_1434_elements(60) & inputPort_2_Daemon_CP_1434_elements(64) & inputPort_2_Daemon_CP_1434_elements(82);
      gj_inputPort_2_Daemon_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81: marked-successors 
    -- CP-element group 81: 	62 
    -- CP-element group 81: 	77 
    -- CP-element group 81: 	58 
    -- CP-element group 81:  members (6) 
      -- CP-element group 81: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_1_479_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_1_479_update_start_
      -- CP-element group 81: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_1_479_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_1_479_Sample/ack
      -- CP-element group 81: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_1_479_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_1_479_Update/req
      -- 
    ack_1663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_1_479_inst_ack_0, ack => inputPort_2_Daemon_CP_1434_elements(81)); -- 
    req_1667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(81), ack => WPIPE_noblock_obuf_2_1_479_inst_req_1); -- 
    -- CP-element group 82:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	102 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	80 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_1_479_Update/ack
      -- CP-element group 82: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_1_479_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_1_479_update_completed_
      -- 
    ack_1668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_1_479_inst_ack_1, ack => inputPort_2_Daemon_CP_1434_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: marked-predecessors 
    -- CP-element group 83: 	87 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_484_update_start_
      -- CP-element group 83: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_484_Update/req
      -- CP-element group 83: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_484_Update/$entry
      -- 
    req_1681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(83), ack => W_data_to_outport_445_delayed_4_0_482_inst_req_1); -- 
    inputPort_2_Daemon_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_2_Daemon_CP_1434_elements(87);
      gj_inputPort_2_Daemon_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	37 
    -- CP-element group 84: successors 
    -- CP-element group 84: marked-successors 
    -- CP-element group 84: 	33 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_484_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_484_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_484_Sample/ack
      -- 
    ack_1677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_445_delayed_4_0_482_inst_ack_0, ack => inputPort_2_Daemon_CP_1434_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_484_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_484_Update/ack
      -- CP-element group 85: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_484_Update/$exit
      -- 
    ack_1682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_445_delayed_4_0_482_inst_ack_1, ack => inputPort_2_Daemon_CP_1434_elements(85)); -- 
    -- CP-element group 86:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: 	68 
    -- CP-element group 86: 	60 
    -- CP-element group 86: marked-predecessors 
    -- CP-element group 86: 	88 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_2_486_Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_2_486_sample_start_
      -- CP-element group 86: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_2_486_Sample/req
      -- 
    req_1690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(86), ack => WPIPE_noblock_obuf_2_2_486_inst_req_0); -- 
    inputPort_2_Daemon_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_1434_elements(85) & inputPort_2_Daemon_CP_1434_elements(68) & inputPort_2_Daemon_CP_1434_elements(60) & inputPort_2_Daemon_CP_1434_elements(88);
      gj_inputPort_2_Daemon_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: marked-successors 
    -- CP-element group 87: 	83 
    -- CP-element group 87: 	66 
    -- CP-element group 87: 	58 
    -- CP-element group 87:  members (6) 
      -- CP-element group 87: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_2_486_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_2_486_update_start_
      -- CP-element group 87: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_2_486_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_2_486_Update/req
      -- CP-element group 87: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_2_486_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_2_486_Sample/ack
      -- 
    ack_1691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_2_486_inst_ack_0, ack => inputPort_2_Daemon_CP_1434_elements(87)); -- 
    req_1695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(87), ack => WPIPE_noblock_obuf_2_2_486_inst_req_1); -- 
    -- CP-element group 88:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	102 
    -- CP-element group 88: marked-successors 
    -- CP-element group 88: 	86 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_2_486_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_2_486_Update/ack
      -- CP-element group 88: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_2_486_Update/$exit
      -- 
    ack_1696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_2_486_inst_ack_1, ack => inputPort_2_Daemon_CP_1434_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	93 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_491_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_491_Update/req
      -- CP-element group 89: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_491_update_start_
      -- 
    req_1709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(89), ack => W_data_to_outport_449_delayed_4_0_489_inst_req_1); -- 
    inputPort_2_Daemon_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_2_Daemon_CP_1434_elements(93);
      gj_inputPort_2_Daemon_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	37 
    -- CP-element group 90: successors 
    -- CP-element group 90: marked-successors 
    -- CP-element group 90: 	33 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_491_Sample/ack
      -- CP-element group 90: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_491_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_491_sample_completed_
      -- 
    ack_1705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_449_delayed_4_0_489_inst_ack_0, ack => inputPort_2_Daemon_CP_1434_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_491_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_491_Update/ack
      -- CP-element group 91: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_491_update_completed_
      -- 
    ack_1710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_449_delayed_4_0_489_inst_ack_1, ack => inputPort_2_Daemon_CP_1434_elements(91)); -- 
    -- CP-element group 92:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: 	72 
    -- CP-element group 92: 	60 
    -- CP-element group 92: marked-predecessors 
    -- CP-element group 92: 	94 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_3_493_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_3_493_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_3_493_Sample/req
      -- 
    req_1718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(92), ack => WPIPE_noblock_obuf_2_3_493_inst_req_0); -- 
    inputPort_2_Daemon_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_1434_elements(91) & inputPort_2_Daemon_CP_1434_elements(72) & inputPort_2_Daemon_CP_1434_elements(60) & inputPort_2_Daemon_CP_1434_elements(94);
      gj_inputPort_2_Daemon_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93: marked-successors 
    -- CP-element group 93: 	89 
    -- CP-element group 93: 	70 
    -- CP-element group 93: 	58 
    -- CP-element group 93:  members (6) 
      -- CP-element group 93: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_3_493_Update/$entry
      -- CP-element group 93: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_3_493_Update/req
      -- CP-element group 93: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_3_493_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_3_493_Sample/ack
      -- CP-element group 93: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_3_493_update_start_
      -- CP-element group 93: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_3_493_Sample/$exit
      -- 
    ack_1719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_3_493_inst_ack_0, ack => inputPort_2_Daemon_CP_1434_elements(93)); -- 
    req_1723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(93), ack => WPIPE_noblock_obuf_2_3_493_inst_req_1); -- 
    -- CP-element group 94:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	102 
    -- CP-element group 94: marked-successors 
    -- CP-element group 94: 	92 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_3_493_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_3_493_Update/ack
      -- CP-element group 94: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_3_493_update_completed_
      -- 
    ack_1724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_3_493_inst_ack_1, ack => inputPort_2_Daemon_CP_1434_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: marked-predecessors 
    -- CP-element group 95: 	99 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_498_update_start_
      -- CP-element group 95: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_498_Update/$entry
      -- CP-element group 95: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_498_Update/req
      -- 
    req_1737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(95), ack => W_data_to_outport_453_delayed_4_0_496_inst_req_1); -- 
    inputPort_2_Daemon_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_2_Daemon_CP_1434_elements(99);
      gj_inputPort_2_Daemon_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	37 
    -- CP-element group 96: successors 
    -- CP-element group 96: marked-successors 
    -- CP-element group 96: 	33 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_498_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_498_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_498_Sample/ack
      -- 
    ack_1733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_453_delayed_4_0_496_inst_ack_0, ack => inputPort_2_Daemon_CP_1434_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_498_Update/ack
      -- CP-element group 97: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_498_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/assign_stmt_498_update_completed_
      -- 
    ack_1738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_453_delayed_4_0_496_inst_ack_1, ack => inputPort_2_Daemon_CP_1434_elements(97)); -- 
    -- CP-element group 98:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: 	60 
    -- CP-element group 98: 	76 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	100 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_4_500_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_4_500_Sample/req
      -- CP-element group 98: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_4_500_sample_start_
      -- 
    req_1746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(98), ack => WPIPE_noblock_obuf_2_4_500_inst_req_0); -- 
    inputPort_2_Daemon_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_1434_elements(97) & inputPort_2_Daemon_CP_1434_elements(60) & inputPort_2_Daemon_CP_1434_elements(76) & inputPort_2_Daemon_CP_1434_elements(100);
      gj_inputPort_2_Daemon_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: marked-successors 
    -- CP-element group 99: 	95 
    -- CP-element group 99: 	74 
    -- CP-element group 99: 	58 
    -- CP-element group 99:  members (6) 
      -- CP-element group 99: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_4_500_Update/$entry
      -- CP-element group 99: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_4_500_Update/req
      -- CP-element group 99: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_4_500_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_4_500_Sample/ack
      -- CP-element group 99: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_4_500_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_4_500_update_start_
      -- 
    ack_1747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_4_500_inst_ack_0, ack => inputPort_2_Daemon_CP_1434_elements(99)); -- 
    req_1751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_1434_elements(99), ack => WPIPE_noblock_obuf_2_4_500_inst_req_1); -- 
    -- CP-element group 100:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100: marked-successors 
    -- CP-element group 100: 	98 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_4_500_Update/ack
      -- CP-element group 100: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_4_500_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/WPIPE_noblock_obuf_2_4_500_update_completed_
      -- 
    ack_1752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_4_500_inst_ack_1, ack => inputPort_2_Daemon_CP_1434_elements(100)); -- 
    -- CP-element group 101:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	9 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	10 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group inputPort_2_Daemon_CP_1434_elements(101) is a control-delay.
    cp_element_101_delay: control_delay_element  generic map(name => " 101_delay", delay_value => 1)  port map(req => inputPort_2_Daemon_CP_1434_elements(9), ack => inputPort_2_Daemon_CP_1434_elements(101), clk => clk, reset =>reset);
    -- CP-element group 102:  join  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	82 
    -- CP-element group 102: 	12 
    -- CP-element group 102: 	13 
    -- CP-element group 102: 	88 
    -- CP-element group 102: 	94 
    -- CP-element group 102: 	100 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	6 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_366/do_while_stmt_367/do_while_stmt_367_loop_body/$exit
      -- 
    inputPort_2_Daemon_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 39) := "inputPort_2_Daemon_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_1434_elements(82) & inputPort_2_Daemon_CP_1434_elements(12) & inputPort_2_Daemon_CP_1434_elements(13) & inputPort_2_Daemon_CP_1434_elements(88) & inputPort_2_Daemon_CP_1434_elements(94) & inputPort_2_Daemon_CP_1434_elements(100);
      gj_inputPort_2_Daemon_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	5 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_366/do_while_stmt_367/loop_exit/$exit
      -- CP-element group 103: 	 branch_block_stmt_366/do_while_stmt_367/loop_exit/ack
      -- 
    ack_1757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_367_branch_ack_0, ack => inputPort_2_Daemon_CP_1434_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	5 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_366/do_while_stmt_367/loop_taken/$exit
      -- CP-element group 104: 	 branch_block_stmt_366/do_while_stmt_367/loop_taken/ack
      -- 
    ack_1761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_367_branch_ack_1, ack => inputPort_2_Daemon_CP_1434_elements(104)); -- 
    -- CP-element group 105:  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	3 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	1 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_366/do_while_stmt_367/$exit
      -- 
    inputPort_2_Daemon_CP_1434_elements(105) <= inputPort_2_Daemon_CP_1434_elements(3);
    inputPort_2_Daemon_do_while_stmt_367_terminator_1762: loop_terminator -- 
      generic map (name => " inputPort_2_Daemon_do_while_stmt_367_terminator_1762", max_iterations_in_flight =>7) 
      port map(loop_body_exit => inputPort_2_Daemon_CP_1434_elements(6),loop_continue => inputPort_2_Daemon_CP_1434_elements(104),loop_terminate => inputPort_2_Daemon_CP_1434_elements(103),loop_back => inputPort_2_Daemon_CP_1434_elements(4),loop_exit => inputPort_2_Daemon_CP_1434_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_369_phi_seq_1508_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_2_Daemon_CP_1434_elements(22);
      inputPort_2_Daemon_CP_1434_elements(25)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_2_Daemon_CP_1434_elements(25);
      inputPort_2_Daemon_CP_1434_elements(26)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_2_Daemon_CP_1434_elements(27);
      inputPort_2_Daemon_CP_1434_elements(23) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_2_Daemon_CP_1434_elements(20);
      inputPort_2_Daemon_CP_1434_elements(29)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_2_Daemon_CP_1434_elements(31);
      inputPort_2_Daemon_CP_1434_elements(30)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_2_Daemon_CP_1434_elements(32);
      inputPort_2_Daemon_CP_1434_elements(21) <= phi_mux_reqs(1);
      phi_stmt_369_phi_seq_1508 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_369_phi_seq_1508") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_2_Daemon_CP_1434_elements(11), 
          phi_sample_ack => inputPort_2_Daemon_CP_1434_elements(18), 
          phi_update_req => inputPort_2_Daemon_CP_1434_elements(14), 
          phi_update_ack => inputPort_2_Daemon_CP_1434_elements(19), 
          phi_mux_ack => inputPort_2_Daemon_CP_1434_elements(24), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_376_phi_seq_1570_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_2_Daemon_CP_1434_elements(46);
      inputPort_2_Daemon_CP_1434_elements(49)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_2_Daemon_CP_1434_elements(49);
      inputPort_2_Daemon_CP_1434_elements(50)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_2_Daemon_CP_1434_elements(51);
      inputPort_2_Daemon_CP_1434_elements(47) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_2_Daemon_CP_1434_elements(44);
      inputPort_2_Daemon_CP_1434_elements(53)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_2_Daemon_CP_1434_elements(55);
      inputPort_2_Daemon_CP_1434_elements(54)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_2_Daemon_CP_1434_elements(56);
      inputPort_2_Daemon_CP_1434_elements(45) <= phi_mux_reqs(1);
      phi_stmt_376_phi_seq_1570 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_376_phi_seq_1570") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_2_Daemon_CP_1434_elements(40), 
          phi_sample_ack => inputPort_2_Daemon_CP_1434_elements(41), 
          phi_update_req => inputPort_2_Daemon_CP_1434_elements(42), 
          phi_update_ack => inputPort_2_Daemon_CP_1434_elements(43), 
          phi_mux_ack => inputPort_2_Daemon_CP_1434_elements(48), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1459_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= inputPort_2_Daemon_CP_1434_elements(7);
        preds(1)  <= inputPort_2_Daemon_CP_1434_elements(8);
        entry_tmerge_1459 : transition_merge -- 
          generic map(name => " entry_tmerge_1459")
          port map (preds => preds, symbol_out => inputPort_2_Daemon_CP_1434_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal EQ_u8_u1_414_414_delayed_4_0_439 : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_421_421_delayed_4_0_449 : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_428_428_delayed_4_0_459 : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_435_435_delayed_4_0_469 : std_logic_vector(0 downto 0);
    signal RPIPE_in_data_2_375_wire : std_logic_vector(31 downto 0);
    signal R_ONE_1_422_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_16_371_wire_constant : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_409_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_412_wire : std_logic_vector(15 downto 0);
    signal SUB_u8_u8_430_wire : std_logic_vector(7 downto 0);
    signal continue_434 : std_logic_vector(0 downto 0);
    signal count_down_369 : std_logic_vector(15 downto 0);
    signal data_to_outport_425 : std_logic_vector(32 downto 0);
    signal data_to_outport_441_delayed_4_0_477 : std_logic_vector(32 downto 0);
    signal data_to_outport_445_delayed_4_0_484 : std_logic_vector(32 downto 0);
    signal data_to_outport_449_delayed_4_0_491 : std_logic_vector(32 downto 0);
    signal data_to_outport_453_delayed_4_0_498 : std_logic_vector(32 downto 0);
    signal dest_id_391 : std_logic_vector(7 downto 0);
    signal input_word_373 : std_logic_vector(31 downto 0);
    signal konst_378_wire_constant : std_logic_vector(7 downto 0);
    signal konst_385_wire_constant : std_logic_vector(15 downto 0);
    signal konst_408_wire_constant : std_logic_vector(15 downto 0);
    signal konst_411_wire_constant : std_logic_vector(15 downto 0);
    signal konst_427_wire_constant : std_logic_vector(7 downto 0);
    signal konst_429_wire_constant : std_logic_vector(7 downto 0);
    signal konst_437_wire_constant : std_logic_vector(7 downto 0);
    signal konst_447_wire_constant : std_logic_vector(7 downto 0);
    signal konst_457_wire_constant : std_logic_vector(7 downto 0);
    signal konst_467_wire_constant : std_logic_vector(7 downto 0);
    signal konst_514_wire_constant : std_logic_vector(0 downto 0);
    signal last_dest_id_376 : std_logic_vector(7 downto 0);
    signal new_packet_387 : std_logic_vector(0 downto 0);
    signal next_count_down_414 : std_logic_vector(15 downto 0);
    signal next_count_down_414_372_buffered : std_logic_vector(15 downto 0);
    signal next_last_dest_id_420 : std_logic_vector(7 downto 0);
    signal next_last_dest_id_420_379_buffered : std_logic_vector(7 downto 0);
    signal pkt_length_395 : std_logic_vector(15 downto 0);
    signal send_to_1_444 : std_logic_vector(0 downto 0);
    signal send_to_2_454 : std_logic_vector(0 downto 0);
    signal send_to_3_464 : std_logic_vector(0 downto 0);
    signal send_to_4_474 : std_logic_vector(0 downto 0);
    signal seq_id_399 : std_logic_vector(7 downto 0);
    signal type_cast_432_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_ONE_1_422_wire_constant <= "1";
    R_ZERO_16_371_wire_constant <= "0000000000000000";
    konst_378_wire_constant <= "00000000";
    konst_385_wire_constant <= "0000000000000000";
    konst_408_wire_constant <= "0000000000000001";
    konst_411_wire_constant <= "0000000000000001";
    konst_427_wire_constant <= "00000001";
    konst_429_wire_constant <= "00000001";
    konst_437_wire_constant <= "00000001";
    konst_447_wire_constant <= "00000010";
    konst_457_wire_constant <= "00000011";
    konst_467_wire_constant <= "00000100";
    konst_514_wire_constant <= "1";
    type_cast_432_wire_constant <= "1";
    phi_stmt_369: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_16_371_wire_constant & next_count_down_414_372_buffered;
      req <= phi_stmt_369_req_0 & phi_stmt_369_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_369",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_369_ack_0,
          idata => idata,
          odata => count_down_369,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_369
    phi_stmt_376: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= konst_378_wire_constant & next_last_dest_id_420_379_buffered;
      req <= phi_stmt_376_req_0 & phi_stmt_376_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_376",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_376_ack_0,
          idata => idata,
          odata => last_dest_id_376,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_376
    -- flow-through select operator MUX_413_inst
    next_count_down_414 <= SUB_u16_u16_409_wire when (new_packet_387(0) /=  '0') else SUB_u16_u16_412_wire;
    -- flow-through select operator MUX_419_inst
    next_last_dest_id_420 <= dest_id_391 when (new_packet_387(0) /=  '0') else last_dest_id_376;
    -- flow-through slice operator slice_390_inst
    dest_id_391 <= input_word_373(31 downto 24);
    -- flow-through slice operator slice_394_inst
    pkt_length_395 <= input_word_373(23 downto 8);
    -- flow-through slice operator slice_398_inst
    seq_id_399 <= input_word_373(7 downto 0);
    W_data_to_outport_441_delayed_4_0_475_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_data_to_outport_441_delayed_4_0_475_inst_req_0;
      W_data_to_outport_441_delayed_4_0_475_inst_ack_0<= wack(0);
      rreq(0) <= W_data_to_outport_441_delayed_4_0_475_inst_req_1;
      W_data_to_outport_441_delayed_4_0_475_inst_ack_1<= rack(0);
      W_data_to_outport_441_delayed_4_0_475_inst : InterlockBuffer generic map ( -- 
        name => "W_data_to_outport_441_delayed_4_0_475_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 33,
        out_data_width => 33,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => data_to_outport_425,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => data_to_outport_441_delayed_4_0_477,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_data_to_outport_445_delayed_4_0_482_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_data_to_outport_445_delayed_4_0_482_inst_req_0;
      W_data_to_outport_445_delayed_4_0_482_inst_ack_0<= wack(0);
      rreq(0) <= W_data_to_outport_445_delayed_4_0_482_inst_req_1;
      W_data_to_outport_445_delayed_4_0_482_inst_ack_1<= rack(0);
      W_data_to_outport_445_delayed_4_0_482_inst : InterlockBuffer generic map ( -- 
        name => "W_data_to_outport_445_delayed_4_0_482_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 33,
        out_data_width => 33,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => data_to_outport_425,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => data_to_outport_445_delayed_4_0_484,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_data_to_outport_449_delayed_4_0_489_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_data_to_outport_449_delayed_4_0_489_inst_req_0;
      W_data_to_outport_449_delayed_4_0_489_inst_ack_0<= wack(0);
      rreq(0) <= W_data_to_outport_449_delayed_4_0_489_inst_req_1;
      W_data_to_outport_449_delayed_4_0_489_inst_ack_1<= rack(0);
      W_data_to_outport_449_delayed_4_0_489_inst : InterlockBuffer generic map ( -- 
        name => "W_data_to_outport_449_delayed_4_0_489_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 33,
        out_data_width => 33,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => data_to_outport_425,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => data_to_outport_449_delayed_4_0_491,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_data_to_outport_453_delayed_4_0_496_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_data_to_outport_453_delayed_4_0_496_inst_req_0;
      W_data_to_outport_453_delayed_4_0_496_inst_ack_0<= wack(0);
      rreq(0) <= W_data_to_outport_453_delayed_4_0_496_inst_req_1;
      W_data_to_outport_453_delayed_4_0_496_inst_ack_1<= rack(0);
      W_data_to_outport_453_delayed_4_0_496_inst : InterlockBuffer generic map ( -- 
        name => "W_data_to_outport_453_delayed_4_0_496_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 33,
        out_data_width => 33,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => data_to_outport_425,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => data_to_outport_453_delayed_4_0_498,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_count_down_414_372_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_count_down_414_372_buf_req_0;
      next_count_down_414_372_buf_ack_0<= wack(0);
      rreq(0) <= next_count_down_414_372_buf_req_1;
      next_count_down_414_372_buf_ack_1<= rack(0);
      next_count_down_414_372_buf : InterlockBuffer generic map ( -- 
        name => "next_count_down_414_372_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_count_down_414,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_count_down_414_372_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_last_dest_id_420_379_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_last_dest_id_420_379_buf_req_0;
      next_last_dest_id_420_379_buf_ack_0<= wack(0);
      rreq(0) <= next_last_dest_id_420_379_buf_req_1;
      next_last_dest_id_420_379_buf_ack_1<= rack(0);
      next_last_dest_id_420_379_buf : InterlockBuffer generic map ( -- 
        name => "next_last_dest_id_420_379_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_last_dest_id_420,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_last_dest_id_420_379_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_373
    process(RPIPE_in_data_2_375_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := RPIPE_in_data_2_375_wire(31 downto 0);
      input_word_373 <= tmp_var; -- 
    end process;
    do_while_stmt_367_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_514_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_367_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_367_branch_req_0,
          ack0 => do_while_stmt_367_branch_ack_0,
          ack1 => do_while_stmt_367_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- flow through binary operator AND_u1_u1_443_inst
    send_to_1_444 <= (EQ_u8_u1_414_414_delayed_4_0_439 and continue_434);
    -- flow through binary operator AND_u1_u1_453_inst
    send_to_2_454 <= (EQ_u8_u1_421_421_delayed_4_0_449 and continue_434);
    -- flow through binary operator AND_u1_u1_463_inst
    send_to_3_464 <= (EQ_u8_u1_428_428_delayed_4_0_459 and continue_434);
    -- flow through binary operator AND_u1_u1_473_inst
    send_to_4_474 <= (EQ_u8_u1_435_435_delayed_4_0_469 and continue_434);
    -- flow through binary operator CONCAT_u1_u33_424_inst
    process(R_ONE_1_422_wire_constant, input_word_373) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ONE_1_422_wire_constant, input_word_373, tmp_var);
      data_to_outport_425 <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u16_u1_386_inst
    process(count_down_369) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(count_down_369, konst_385_wire_constant, tmp_var);
      new_packet_387 <= tmp_var; --
    end process;
    -- shared split operator group (6) : EQ_u8_u1_438_inst 
    ApIntEq_group_6: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 4);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= next_last_dest_id_420;
      EQ_u8_u1_414_414_delayed_4_0_439 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u8_u1_438_inst_req_0;
      EQ_u8_u1_438_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u8_u1_438_inst_req_1;
      EQ_u8_u1_438_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_6_gI: SplitGuardInterface generic map(name => "ApIntEq_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000001",
          constant_width => 8,
          buffering  => 4,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : EQ_u8_u1_448_inst 
    ApIntEq_group_7: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 4);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= next_last_dest_id_420;
      EQ_u8_u1_421_421_delayed_4_0_449 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u8_u1_448_inst_req_0;
      EQ_u8_u1_448_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u8_u1_448_inst_req_1;
      EQ_u8_u1_448_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_7_gI: SplitGuardInterface generic map(name => "ApIntEq_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000010",
          constant_width => 8,
          buffering  => 4,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : EQ_u8_u1_458_inst 
    ApIntEq_group_8: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 4);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= next_last_dest_id_420;
      EQ_u8_u1_428_428_delayed_4_0_459 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u8_u1_458_inst_req_0;
      EQ_u8_u1_458_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u8_u1_458_inst_req_1;
      EQ_u8_u1_458_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_8_gI: SplitGuardInterface generic map(name => "ApIntEq_group_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_8",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000011",
          constant_width => 8,
          buffering  => 4,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : EQ_u8_u1_468_inst 
    ApIntEq_group_9: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 4);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= next_last_dest_id_420;
      EQ_u8_u1_435_435_delayed_4_0_469 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u8_u1_468_inst_req_0;
      EQ_u8_u1_468_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u8_u1_468_inst_req_1;
      EQ_u8_u1_468_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_9_gI: SplitGuardInterface generic map(name => "ApIntEq_group_9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_9",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000100",
          constant_width => 8,
          buffering  => 4,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- flow through binary operator SUB_u16_u16_409_inst
    SUB_u16_u16_409_wire <= std_logic_vector(unsigned(pkt_length_395) - unsigned(konst_408_wire_constant));
    -- flow through binary operator SUB_u16_u16_412_inst
    SUB_u16_u16_412_wire <= std_logic_vector(unsigned(count_down_369) - unsigned(konst_411_wire_constant));
    -- flow through binary operator SUB_u8_u8_430_inst
    SUB_u8_u8_430_wire <= std_logic_vector(unsigned(next_last_dest_id_420) - unsigned(konst_429_wire_constant));
    -- shared inport operator group (0) : RPIPE_in_data_2_375_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_in_data_2_375_inst_req_0;
      RPIPE_in_data_2_375_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_in_data_2_375_inst_req_1;
      RPIPE_in_data_2_375_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_in_data_2_375_wire <= data_out(31 downto 0);
      in_data_2_read_0_gI: SplitGuardInterface generic map(name => "in_data_2_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      in_data_2_read_0: InputPortRevised -- 
        generic map ( name => "in_data_2_read_0", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => in_data_2_pipe_read_req(0),
          oack => in_data_2_pipe_read_ack(0),
          odata => in_data_2_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_noblock_obuf_2_1_479_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_2_1_479_inst_req_0;
      WPIPE_noblock_obuf_2_1_479_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_2_1_479_inst_req_1;
      WPIPE_noblock_obuf_2_1_479_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_1_444(0);
      data_in <= data_to_outport_441_delayed_4_0_477;
      noblock_obuf_2_1_write_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_1_write_0: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_2_1", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_2_1_pipe_write_req(0),
          oack => noblock_obuf_2_1_pipe_write_ack(0),
          odata => noblock_obuf_2_1_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_noblock_obuf_2_2_486_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_2_2_486_inst_req_0;
      WPIPE_noblock_obuf_2_2_486_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_2_2_486_inst_req_1;
      WPIPE_noblock_obuf_2_2_486_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_2_454(0);
      data_in <= data_to_outport_445_delayed_4_0_484;
      noblock_obuf_2_2_write_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_2_write_1: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_2_2", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_2_2_pipe_write_req(0),
          oack => noblock_obuf_2_2_pipe_write_ack(0),
          odata => noblock_obuf_2_2_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_noblock_obuf_2_3_493_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_2_3_493_inst_req_0;
      WPIPE_noblock_obuf_2_3_493_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_2_3_493_inst_req_1;
      WPIPE_noblock_obuf_2_3_493_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_3_464(0);
      data_in <= data_to_outport_449_delayed_4_0_491;
      noblock_obuf_2_3_write_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_3_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_3_write_2: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_2_3", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_2_3_pipe_write_req(0),
          oack => noblock_obuf_2_3_pipe_write_ack(0),
          odata => noblock_obuf_2_3_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_noblock_obuf_2_4_500_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_2_4_500_inst_req_0;
      WPIPE_noblock_obuf_2_4_500_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_2_4_500_inst_req_1;
      WPIPE_noblock_obuf_2_4_500_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_4_474(0);
      data_in <= data_to_outport_453_delayed_4_0_498;
      noblock_obuf_2_4_write_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_4_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_4_write_3: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_2_4", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_2_4_pipe_write_req(0),
          oack => noblock_obuf_2_4_pipe_write_ack(0),
          odata => noblock_obuf_2_4_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared call operator group (0) : call_updateCounter_expr_433_inst 
    updateCounter_call_group_0: Block -- 
      signal data_in: std_logic_vector(16 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_updateCounter_expr_433_inst_req_0;
      call_updateCounter_expr_433_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_updateCounter_expr_433_inst_req_1;
      call_updateCounter_expr_433_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      updateCounter_call_group_0_gI: SplitGuardInterface generic map(name => "updateCounter_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_427_wire_constant & SUB_u8_u8_430_wire & type_cast_432_wire_constant;
      continue_434 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 17,
        owidth => 17,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => updateCounter_call_reqs(0),
          ackR => updateCounter_call_acks(0),
          dataR => updateCounter_call_data(16 downto 0),
          tagR => updateCounter_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => updateCounter_return_acks(0), -- cross-over
          ackL => updateCounter_return_reqs(0), -- cross-over
          dataL => updateCounter_return_data(0 downto 0),
          tagL => updateCounter_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end inputPort_2_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity inputPort_3_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    in_data_3_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_3_pipe_read_data : in   std_logic_vector(31 downto 0);
    noblock_obuf_3_2_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_2_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_3_3_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_3_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_3_4_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_4_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_3_1_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_1_pipe_write_data : out  std_logic_vector(32 downto 0);
    updateCounter_call_reqs : out  std_logic_vector(0 downto 0);
    updateCounter_call_acks : in   std_logic_vector(0 downto 0);
    updateCounter_call_data : out  std_logic_vector(16 downto 0);
    updateCounter_call_tag  :  out  std_logic_vector(0 downto 0);
    updateCounter_return_reqs : out  std_logic_vector(0 downto 0);
    updateCounter_return_acks : in   std_logic_vector(0 downto 0);
    updateCounter_return_data : in   std_logic_vector(0 downto 0);
    updateCounter_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity inputPort_3_Daemon;
architecture inputPort_3_Daemon_arch of inputPort_3_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal inputPort_3_Daemon_CP_1763_start: Boolean;
  signal inputPort_3_Daemon_CP_1763_symbol: Boolean;
  -- volatile/operator module components. 
  component updateCounter is -- 
    generic (tag_length : integer); 
    port ( -- 
      input_port : in  std_logic_vector(7 downto 0);
      output_port : in  std_logic_vector(7 downto 0);
      up : in  std_logic_vector(0 downto 0);
      continue : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(3 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(1 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(1 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal WPIPE_noblock_obuf_3_4_652_inst_ack_1 : boolean;
  signal W_data_to_outport_569_delayed_4_0_627_inst_ack_1 : boolean;
  signal W_data_to_outport_581_delayed_4_0_648_inst_ack_1 : boolean;
  signal W_data_to_outport_573_delayed_4_0_634_inst_ack_0 : boolean;
  signal W_data_to_outport_569_delayed_4_0_627_inst_req_1 : boolean;
  signal EQ_u8_u1_620_inst_ack_0 : boolean;
  signal W_data_to_outport_577_delayed_4_0_641_inst_ack_0 : boolean;
  signal EQ_u8_u1_620_inst_req_1 : boolean;
  signal W_data_to_outport_577_delayed_4_0_641_inst_req_0 : boolean;
  signal EQ_u8_u1_600_inst_ack_0 : boolean;
  signal next_last_dest_id_572_531_buf_req_0 : boolean;
  signal WPIPE_noblock_obuf_3_1_631_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_3_3_645_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_3_3_645_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_3_1_631_inst_ack_0 : boolean;
  signal call_updateCounter_expr_585_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_3_4_652_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_3_1_631_inst_ack_1 : boolean;
  signal W_data_to_outport_573_delayed_4_0_634_inst_req_0 : boolean;
  signal EQ_u8_u1_610_inst_ack_0 : boolean;
  signal EQ_u8_u1_610_inst_req_0 : boolean;
  signal next_last_dest_id_572_531_buf_ack_1 : boolean;
  signal WPIPE_noblock_obuf_3_4_652_inst_req_0 : boolean;
  signal next_last_dest_id_572_531_buf_req_1 : boolean;
  signal WPIPE_noblock_obuf_3_2_638_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_3_4_652_inst_req_1 : boolean;
  signal next_last_dest_id_572_531_buf_ack_0 : boolean;
  signal W_data_to_outport_581_delayed_4_0_648_inst_req_1 : boolean;
  signal do_while_stmt_519_branch_ack_0 : boolean;
  signal EQ_u8_u1_610_inst_ack_1 : boolean;
  signal EQ_u8_u1_600_inst_req_0 : boolean;
  signal EQ_u8_u1_620_inst_ack_1 : boolean;
  signal EQ_u8_u1_590_inst_ack_0 : boolean;
  signal EQ_u8_u1_590_inst_req_0 : boolean;
  signal EQ_u8_u1_620_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_3_2_638_inst_req_1 : boolean;
  signal EQ_u8_u1_590_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_3_1_631_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_3_3_645_inst_req_1 : boolean;
  signal call_updateCounter_expr_585_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_3_3_645_inst_req_0 : boolean;
  signal W_data_to_outport_569_delayed_4_0_627_inst_ack_0 : boolean;
  signal EQ_u8_u1_610_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_3_2_638_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_3_2_638_inst_ack_0 : boolean;
  signal EQ_u8_u1_590_inst_ack_1 : boolean;
  signal phi_stmt_528_ack_0 : boolean;
  signal W_data_to_outport_569_delayed_4_0_627_inst_req_0 : boolean;
  signal call_updateCounter_expr_585_inst_ack_0 : boolean;
  signal W_data_to_outport_581_delayed_4_0_648_inst_ack_0 : boolean;
  signal call_updateCounter_expr_585_inst_req_0 : boolean;
  signal W_data_to_outport_577_delayed_4_0_641_inst_ack_1 : boolean;
  signal W_data_to_outport_577_delayed_4_0_641_inst_req_1 : boolean;
  signal W_data_to_outport_573_delayed_4_0_634_inst_ack_1 : boolean;
  signal W_data_to_outport_581_delayed_4_0_648_inst_req_0 : boolean;
  signal phi_stmt_528_req_0 : boolean;
  signal do_while_stmt_519_branch_ack_1 : boolean;
  signal EQ_u8_u1_600_inst_ack_1 : boolean;
  signal W_data_to_outport_573_delayed_4_0_634_inst_req_1 : boolean;
  signal EQ_u8_u1_600_inst_req_1 : boolean;
  signal do_while_stmt_519_branch_req_0 : boolean;
  signal phi_stmt_521_req_1 : boolean;
  signal phi_stmt_521_req_0 : boolean;
  signal phi_stmt_521_ack_0 : boolean;
  signal next_count_down_566_524_buf_req_0 : boolean;
  signal next_count_down_566_524_buf_ack_0 : boolean;
  signal next_count_down_566_524_buf_req_1 : boolean;
  signal next_count_down_566_524_buf_ack_1 : boolean;
  signal RPIPE_in_data_3_527_inst_req_0 : boolean;
  signal RPIPE_in_data_3_527_inst_ack_0 : boolean;
  signal RPIPE_in_data_3_527_inst_req_1 : boolean;
  signal RPIPE_in_data_3_527_inst_ack_1 : boolean;
  signal phi_stmt_528_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "inputPort_3_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  inputPort_3_Daemon_CP_1763_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "inputPort_3_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_3_Daemon_CP_1763_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= inputPort_3_Daemon_CP_1763_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_3_Daemon_CP_1763_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  inputPort_3_Daemon_CP_1763: Block -- control-path 
    signal inputPort_3_Daemon_CP_1763_elements: BooleanArray(105 downto 0);
    -- 
  begin -- 
    inputPort_3_Daemon_CP_1763_elements(0) <= inputPort_3_Daemon_CP_1763_start;
    inputPort_3_Daemon_CP_1763_symbol <= inputPort_3_Daemon_CP_1763_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_518/$entry
      -- CP-element group 0: 	 branch_block_stmt_518/branch_block_stmt_518__entry__
      -- CP-element group 0: 	 branch_block_stmt_518/do_while_stmt_519__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	105 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_518/$exit
      -- CP-element group 1: 	 branch_block_stmt_518/branch_block_stmt_518__exit__
      -- CP-element group 1: 	 branch_block_stmt_518/do_while_stmt_519__exit__
      -- 
    inputPort_3_Daemon_CP_1763_elements(1) <= inputPort_3_Daemon_CP_1763_elements(105);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_518/do_while_stmt_519/$entry
      -- CP-element group 2: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519__entry__
      -- 
    inputPort_3_Daemon_CP_1763_elements(2) <= inputPort_3_Daemon_CP_1763_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	105 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519__exit__
      -- 
    -- Element group inputPort_3_Daemon_CP_1763_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_518/do_while_stmt_519/loop_back
      -- 
    -- Element group inputPort_3_Daemon_CP_1763_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	103 
    -- CP-element group 5: 	104 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_518/do_while_stmt_519/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_518/do_while_stmt_519/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_518/do_while_stmt_519/condition_done
      -- 
    inputPort_3_Daemon_CP_1763_elements(5) <= inputPort_3_Daemon_CP_1763_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	102 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_518/do_while_stmt_519/loop_body_done
      -- 
    inputPort_3_Daemon_CP_1763_elements(6) <= inputPort_3_Daemon_CP_1763_elements(102);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	20 
    -- CP-element group 7: 	44 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/back_edge_to_loop_body
      -- 
    inputPort_3_Daemon_CP_1763_elements(7) <= inputPort_3_Daemon_CP_1763_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	22 
    -- CP-element group 8: 	46 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/first_time_through_loop_body
      -- 
    inputPort_3_Daemon_CP_1763_elements(8) <= inputPort_3_Daemon_CP_1763_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	101 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	17 
    -- CP-element group 9: 	33 
    -- CP-element group 9: 	38 
    -- CP-element group 9: 	39 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_525_sample_start_
      -- 
    -- Element group inputPort_3_Daemon_CP_1763_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	101 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/condition_evaluated
      -- 
    condition_evaluated_1787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(10), ack => do_while_stmt_519_branch_req_0); -- 
    inputPort_3_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_1763_elements(101) & inputPort_3_Daemon_CP_1763_elements(15);
      gj_inputPort_3_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	16 
    -- CP-element group 11: 	38 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	40 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_521_sample_start__ps
      -- 
    inputPort_3_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_1763_elements(9) & inputPort_3_Daemon_CP_1763_elements(16) & inputPort_3_Daemon_CP_1763_elements(38) & inputPort_3_Daemon_CP_1763_elements(15);
      gj_inputPort_3_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	18 
    -- CP-element group 12: 	36 
    -- CP-element group 12: 	41 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	102 
    -- CP-element group 12: 	13 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	16 
    -- CP-element group 12: 	38 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_521_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_525_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_528_sample_completed_
      -- 
    inputPort_3_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_1763_elements(18) & inputPort_3_Daemon_CP_1763_elements(36) & inputPort_3_Daemon_CP_1763_elements(41);
      gj_inputPort_3_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	102 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/aggregated_phi_sample_ack_d
      -- 
    -- Element group inputPort_3_Daemon_CP_1763_elements(13) is a control-delay.
    cp_element_13_delay: control_delay_element  generic map(name => " 13_delay", delay_value => 1)  port map(req => inputPort_3_Daemon_CP_1763_elements(12), ack => inputPort_3_Daemon_CP_1763_elements(13), clk => clk, reset =>reset);
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	17 
    -- CP-element group 14: 	33 
    -- CP-element group 14: 	39 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	35 
    -- CP-element group 14: 	42 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/aggregated_phi_update_req
      -- CP-element group 14: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_521_update_start__ps
      -- 
    inputPort_3_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_1763_elements(17) & inputPort_3_Daemon_CP_1763_elements(33) & inputPort_3_Daemon_CP_1763_elements(39);
      gj_inputPort_3_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	19 
    -- CP-element group 15: 	37 
    -- CP-element group 15: 	43 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/aggregated_phi_update_ack
      -- 
    inputPort_3_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_1763_elements(19) & inputPort_3_Daemon_CP_1763_elements(37) & inputPort_3_Daemon_CP_1763_elements(43);
      gj_inputPort_3_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	11 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_521_sample_start_
      -- 
    inputPort_3_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_1763_elements(9) & inputPort_3_Daemon_CP_1763_elements(12);
      gj_inputPort_3_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	9 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	59 
    -- CP-element group 17: 	67 
    -- CP-element group 17: 	71 
    -- CP-element group 17: 	75 
    -- CP-element group 17: 	63 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	14 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_521_update_start_
      -- 
    inputPort_3_Daemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_1763_elements(9) & inputPort_3_Daemon_CP_1763_elements(59) & inputPort_3_Daemon_CP_1763_elements(67) & inputPort_3_Daemon_CP_1763_elements(71) & inputPort_3_Daemon_CP_1763_elements(75) & inputPort_3_Daemon_CP_1763_elements(63);
      gj_inputPort_3_Daemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_521_sample_completed__ps
      -- 
    -- Element group inputPort_3_Daemon_CP_1763_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	57 
    -- CP-element group 19: 	15 
    -- CP-element group 19: 	65 
    -- CP-element group 19: 	61 
    -- CP-element group 19: 	69 
    -- CP-element group 19: 	73 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_521_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_521_update_completed__ps
      -- 
    -- Element group inputPort_3_Daemon_CP_1763_elements(19) is bound as output of CP function.
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	7 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_521_loopback_trigger
      -- 
    inputPort_3_Daemon_CP_1763_elements(20) <= inputPort_3_Daemon_CP_1763_elements(7);
    -- CP-element group 21:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_521_loopback_sample_req
      -- CP-element group 21: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_521_loopback_sample_req_ps
      -- 
    phi_stmt_521_loopback_sample_req_1803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_521_loopback_sample_req_1803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(21), ack => phi_stmt_521_req_1); -- 
    -- Element group inputPort_3_Daemon_CP_1763_elements(21) is bound as output of CP function.
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	8 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_521_entry_trigger
      -- 
    inputPort_3_Daemon_CP_1763_elements(22) <= inputPort_3_Daemon_CP_1763_elements(8);
    -- CP-element group 23:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_521_entry_sample_req
      -- CP-element group 23: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_521_entry_sample_req_ps
      -- 
    phi_stmt_521_entry_sample_req_1806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_521_entry_sample_req_1806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(23), ack => phi_stmt_521_req_0); -- 
    -- Element group inputPort_3_Daemon_CP_1763_elements(23) is bound as output of CP function.
    -- CP-element group 24:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_521_phi_mux_ack
      -- CP-element group 24: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_521_phi_mux_ack_ps
      -- 
    phi_stmt_521_phi_mux_ack_1809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_521_ack_0, ack => inputPort_3_Daemon_CP_1763_elements(24)); -- 
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_ZERO_16_523_sample_start__ps
      -- CP-element group 25: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_ZERO_16_523_sample_completed__ps
      -- CP-element group 25: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_ZERO_16_523_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_ZERO_16_523_sample_completed_
      -- 
    -- Element group inputPort_3_Daemon_CP_1763_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_ZERO_16_523_update_start__ps
      -- CP-element group 26: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_ZERO_16_523_update_start_
      -- 
    -- Element group inputPort_3_Daemon_CP_1763_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	28 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_ZERO_16_523_update_completed__ps
      -- 
    inputPort_3_Daemon_CP_1763_elements(27) <= inputPort_3_Daemon_CP_1763_elements(28);
    -- CP-element group 28:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	27 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_ZERO_16_523_update_completed_
      -- 
    -- Element group inputPort_3_Daemon_CP_1763_elements(28) is a control-delay.
    cp_element_28_delay: control_delay_element  generic map(name => " 28_delay", delay_value => 1)  port map(req => inputPort_3_Daemon_CP_1763_elements(26), ack => inputPort_3_Daemon_CP_1763_elements(28), clk => clk, reset =>reset);
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_count_down_524_sample_start__ps
      -- CP-element group 29: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_count_down_524_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_count_down_524_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_count_down_524_Sample/req
      -- 
    req_1830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(29), ack => next_count_down_566_524_buf_req_0); -- 
    -- Element group inputPort_3_Daemon_CP_1763_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_count_down_524_update_start__ps
      -- CP-element group 30: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_count_down_524_update_start_
      -- CP-element group 30: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_count_down_524_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_count_down_524_Update/req
      -- 
    req_1835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(30), ack => next_count_down_566_524_buf_req_1); -- 
    -- Element group inputPort_3_Daemon_CP_1763_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_count_down_524_sample_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_count_down_524_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_count_down_524_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_count_down_524_Sample/ack
      -- 
    ack_1831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_566_524_buf_ack_0, ack => inputPort_3_Daemon_CP_1763_elements(31)); -- 
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_count_down_524_update_completed__ps
      -- CP-element group 32: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_count_down_524_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_count_down_524_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_count_down_524_Update/ack
      -- 
    ack_1836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_566_524_buf_ack_1, ack => inputPort_3_Daemon_CP_1763_elements(32)); -- 
    -- CP-element group 33:  join  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	9 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	59 
    -- CP-element group 33: 	96 
    -- CP-element group 33: 	67 
    -- CP-element group 33: 	90 
    -- CP-element group 33: 	84 
    -- CP-element group 33: 	78 
    -- CP-element group 33: 	71 
    -- CP-element group 33: 	75 
    -- CP-element group 33: 	63 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	14 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_525_update_start_
      -- 
    inputPort_3_Daemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_1763_elements(9) & inputPort_3_Daemon_CP_1763_elements(59) & inputPort_3_Daemon_CP_1763_elements(96) & inputPort_3_Daemon_CP_1763_elements(67) & inputPort_3_Daemon_CP_1763_elements(90) & inputPort_3_Daemon_CP_1763_elements(84) & inputPort_3_Daemon_CP_1763_elements(78) & inputPort_3_Daemon_CP_1763_elements(71) & inputPort_3_Daemon_CP_1763_elements(75) & inputPort_3_Daemon_CP_1763_elements(63);
      gj_inputPort_3_Daemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	11 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	37 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/RPIPE_in_data_3_527_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/RPIPE_in_data_3_527_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/RPIPE_in_data_3_527_Sample/rr
      -- 
    rr_1849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(34), ack => RPIPE_in_data_3_527_inst_req_0); -- 
    inputPort_3_Daemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_1763_elements(11) & inputPort_3_Daemon_CP_1763_elements(37);
      gj_inputPort_3_Daemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	14 
    -- CP-element group 35: 	36 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/RPIPE_in_data_3_527_update_start_
      -- CP-element group 35: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/RPIPE_in_data_3_527_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/RPIPE_in_data_3_527_Update/cr
      -- 
    cr_1854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(35), ack => RPIPE_in_data_3_527_inst_req_1); -- 
    inputPort_3_Daemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_1763_elements(14) & inputPort_3_Daemon_CP_1763_elements(36);
      gj_inputPort_3_Daemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	12 
    -- CP-element group 36: 	35 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/RPIPE_in_data_3_527_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/RPIPE_in_data_3_527_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/RPIPE_in_data_3_527_Sample/ra
      -- 
    ra_1850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_3_527_inst_ack_0, ack => inputPort_3_Daemon_CP_1763_elements(36)); -- 
    -- CP-element group 37:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	96 
    -- CP-element group 37: 	57 
    -- CP-element group 37: 	15 
    -- CP-element group 37: 	65 
    -- CP-element group 37: 	90 
    -- CP-element group 37: 	61 
    -- CP-element group 37: 	84 
    -- CP-element group 37: 	78 
    -- CP-element group 37: 	69 
    -- CP-element group 37: 	73 
    -- CP-element group 37: marked-successors 
    -- CP-element group 37: 	34 
    -- CP-element group 37:  members (16) 
      -- CP-element group 37: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_643_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_650_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_629_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_643_Sample/req
      -- CP-element group 37: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_650_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_636_Sample/req
      -- CP-element group 37: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_636_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_643_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_636_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_629_Sample/req
      -- CP-element group 37: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_650_Sample/req
      -- CP-element group 37: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_629_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_525_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/RPIPE_in_data_3_527_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/RPIPE_in_data_3_527_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/RPIPE_in_data_3_527_Update/ca
      -- 
    ca_1855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_3_527_inst_ack_1, ack => inputPort_3_Daemon_CP_1763_elements(37)); -- 
    req_2061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(37), ack => W_data_to_outport_581_delayed_4_0_648_inst_req_0); -- 
    req_2033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(37), ack => W_data_to_outport_577_delayed_4_0_641_inst_req_0); -- 
    req_2005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(37), ack => W_data_to_outport_573_delayed_4_0_634_inst_req_0); -- 
    req_1977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(37), ack => W_data_to_outport_569_delayed_4_0_627_inst_req_0); -- 
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	9 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	12 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	11 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_528_sample_start_
      -- 
    inputPort_3_Daemon_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_1763_elements(9) & inputPort_3_Daemon_CP_1763_elements(12);
      gj_inputPort_3_Daemon_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  join  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	9 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	59 
    -- CP-element group 39: 	67 
    -- CP-element group 39: 	71 
    -- CP-element group 39: 	75 
    -- CP-element group 39: 	63 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	14 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_528_update_start_
      -- 
    inputPort_3_Daemon_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_1763_elements(9) & inputPort_3_Daemon_CP_1763_elements(59) & inputPort_3_Daemon_CP_1763_elements(67) & inputPort_3_Daemon_CP_1763_elements(71) & inputPort_3_Daemon_CP_1763_elements(75) & inputPort_3_Daemon_CP_1763_elements(63);
      gj_inputPort_3_Daemon_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	11 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_528_sample_start__ps
      -- 
    inputPort_3_Daemon_CP_1763_elements(40) <= inputPort_3_Daemon_CP_1763_elements(11);
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	12 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_528_sample_completed__ps
      -- 
    -- Element group inputPort_3_Daemon_CP_1763_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	14 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_528_update_start__ps
      -- 
    inputPort_3_Daemon_CP_1763_elements(42) <= inputPort_3_Daemon_CP_1763_elements(14);
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	57 
    -- CP-element group 43: 	15 
    -- CP-element group 43: 	65 
    -- CP-element group 43: 	61 
    -- CP-element group 43: 	69 
    -- CP-element group 43: 	73 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_528_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_528_update_completed__ps
      -- 
    -- Element group inputPort_3_Daemon_CP_1763_elements(43) is bound as output of CP function.
    -- CP-element group 44:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	7 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_528_loopback_trigger
      -- 
    inputPort_3_Daemon_CP_1763_elements(44) <= inputPort_3_Daemon_CP_1763_elements(7);
    -- CP-element group 45:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_528_loopback_sample_req
      -- CP-element group 45: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_528_loopback_sample_req_ps
      -- 
    phi_stmt_528_loopback_sample_req_1865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_528_loopback_sample_req_1865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(45), ack => phi_stmt_528_req_1); -- 
    -- Element group inputPort_3_Daemon_CP_1763_elements(45) is bound as output of CP function.
    -- CP-element group 46:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	8 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_528_entry_trigger
      -- 
    inputPort_3_Daemon_CP_1763_elements(46) <= inputPort_3_Daemon_CP_1763_elements(8);
    -- CP-element group 47:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_528_entry_sample_req_ps
      -- CP-element group 47: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_528_entry_sample_req
      -- 
    phi_stmt_528_entry_sample_req_1868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_528_entry_sample_req_1868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(47), ack => phi_stmt_528_req_0); -- 
    -- Element group inputPort_3_Daemon_CP_1763_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_528_phi_mux_ack_ps
      -- CP-element group 48: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/phi_stmt_528_phi_mux_ack
      -- 
    phi_stmt_528_phi_mux_ack_1871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_528_ack_0, ack => inputPort_3_Daemon_CP_1763_elements(48)); -- 
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/konst_530_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/konst_530_sample_completed__ps
      -- CP-element group 49: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/konst_530_sample_start__ps
      -- CP-element group 49: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/konst_530_sample_start_
      -- 
    -- Element group inputPort_3_Daemon_CP_1763_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (2) 
      -- CP-element group 50: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/konst_530_update_start_
      -- CP-element group 50: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/konst_530_update_start__ps
      -- 
    -- Element group inputPort_3_Daemon_CP_1763_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	52 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/konst_530_update_completed__ps
      -- 
    inputPort_3_Daemon_CP_1763_elements(51) <= inputPort_3_Daemon_CP_1763_elements(52);
    -- CP-element group 52:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	51 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/konst_530_update_completed_
      -- 
    -- Element group inputPort_3_Daemon_CP_1763_elements(52) is a control-delay.
    cp_element_52_delay: control_delay_element  generic map(name => " 52_delay", delay_value => 1)  port map(req => inputPort_3_Daemon_CP_1763_elements(50), ack => inputPort_3_Daemon_CP_1763_elements(52), clk => clk, reset =>reset);
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_last_dest_id_531_sample_start__ps
      -- CP-element group 53: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_last_dest_id_531_Sample/req
      -- CP-element group 53: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_last_dest_id_531_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_last_dest_id_531_Sample/$entry
      -- 
    req_1892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(53), ack => next_last_dest_id_572_531_buf_req_0); -- 
    -- Element group inputPort_3_Daemon_CP_1763_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_last_dest_id_531_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_last_dest_id_531_update_start__ps
      -- CP-element group 54: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_last_dest_id_531_Update/req
      -- CP-element group 54: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_last_dest_id_531_update_start_
      -- 
    req_1897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(54), ack => next_last_dest_id_572_531_buf_req_1); -- 
    -- Element group inputPort_3_Daemon_CP_1763_elements(54) is bound as output of CP function.
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_last_dest_id_531_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_last_dest_id_531_Sample/ack
      -- CP-element group 55: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_last_dest_id_531_sample_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_last_dest_id_531_sample_completed_
      -- 
    ack_1893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_572_531_buf_ack_0, ack => inputPort_3_Daemon_CP_1763_elements(55)); -- 
    -- CP-element group 56:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_last_dest_id_531_update_completed__ps
      -- CP-element group 56: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_last_dest_id_531_Update/ack
      -- CP-element group 56: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_last_dest_id_531_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/R_next_last_dest_id_531_update_completed_
      -- 
    ack_1898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_572_531_buf_ack_1, ack => inputPort_3_Daemon_CP_1763_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	19 
    -- CP-element group 57: 	37 
    -- CP-element group 57: 	43 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/call_updateCounter_expr_585_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/call_updateCounter_expr_585_Sample/req
      -- CP-element group 57: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/call_updateCounter_expr_585_Sample/$entry
      -- 
    req_1907_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1907_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(57), ack => call_updateCounter_expr_585_inst_req_0); -- 
    inputPort_3_Daemon_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_1763_elements(19) & inputPort_3_Daemon_CP_1763_elements(37) & inputPort_3_Daemon_CP_1763_elements(43);
      gj_inputPort_3_Daemon_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	87 
    -- CP-element group 58: 	99 
    -- CP-element group 58: 	93 
    -- CP-element group 58: 	81 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/call_updateCounter_expr_585_Update/req
      -- CP-element group 58: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/call_updateCounter_expr_585_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/call_updateCounter_expr_585_update_start_
      -- 
    req_1912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(58), ack => call_updateCounter_expr_585_inst_req_1); -- 
    inputPort_3_Daemon_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_1763_elements(87) & inputPort_3_Daemon_CP_1763_elements(99) & inputPort_3_Daemon_CP_1763_elements(93) & inputPort_3_Daemon_CP_1763_elements(81);
      gj_inputPort_3_Daemon_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: marked-successors 
    -- CP-element group 59: 	17 
    -- CP-element group 59: 	33 
    -- CP-element group 59: 	39 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/call_updateCounter_expr_585_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/call_updateCounter_expr_585_Sample/ack
      -- CP-element group 59: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/call_updateCounter_expr_585_Sample/$exit
      -- 
    ack_1908_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_updateCounter_expr_585_inst_ack_0, ack => inputPort_3_Daemon_CP_1763_elements(59)); -- 
    -- CP-element group 60:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	86 
    -- CP-element group 60: 	98 
    -- CP-element group 60: 	92 
    -- CP-element group 60: 	80 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/call_updateCounter_expr_585_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/call_updateCounter_expr_585_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/call_updateCounter_expr_585_update_completed_
      -- 
    ack_1913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_updateCounter_expr_585_inst_ack_1, ack => inputPort_3_Daemon_CP_1763_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	19 
    -- CP-element group 61: 	37 
    -- CP-element group 61: 	43 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_590_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_590_Sample/rr
      -- CP-element group 61: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_590_sample_start_
      -- 
    rr_1921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(61), ack => EQ_u8_u1_590_inst_req_0); -- 
    inputPort_3_Daemon_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_1763_elements(19) & inputPort_3_Daemon_CP_1763_elements(37) & inputPort_3_Daemon_CP_1763_elements(43);
      gj_inputPort_3_Daemon_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	81 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_590_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_590_update_start_
      -- CP-element group 62: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_590_Update/cr
      -- 
    cr_1926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(62), ack => EQ_u8_u1_590_inst_req_1); -- 
    inputPort_3_Daemon_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_3_Daemon_CP_1763_elements(81);
      gj_inputPort_3_Daemon_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	17 
    -- CP-element group 63: 	33 
    -- CP-element group 63: 	39 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_590_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_590_Sample/ra
      -- CP-element group 63: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_590_Sample/$exit
      -- 
    ra_1922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_590_inst_ack_0, ack => inputPort_3_Daemon_CP_1763_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	80 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_590_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_590_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_590_Update/ca
      -- 
    ca_1927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_590_inst_ack_1, ack => inputPort_3_Daemon_CP_1763_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	19 
    -- CP-element group 65: 	37 
    -- CP-element group 65: 	43 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_600_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_600_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_600_Sample/rr
      -- 
    rr_1935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(65), ack => EQ_u8_u1_600_inst_req_0); -- 
    inputPort_3_Daemon_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_1763_elements(19) & inputPort_3_Daemon_CP_1763_elements(37) & inputPort_3_Daemon_CP_1763_elements(43);
      gj_inputPort_3_Daemon_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	87 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_600_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_600_update_start_
      -- CP-element group 66: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_600_Update/cr
      -- 
    cr_1940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(66), ack => EQ_u8_u1_600_inst_req_1); -- 
    inputPort_3_Daemon_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_3_Daemon_CP_1763_elements(87);
      gj_inputPort_3_Daemon_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	17 
    -- CP-element group 67: 	33 
    -- CP-element group 67: 	39 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_600_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_600_Sample/ra
      -- CP-element group 67: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_600_sample_completed_
      -- 
    ra_1936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_600_inst_ack_0, ack => inputPort_3_Daemon_CP_1763_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	86 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_600_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_600_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_600_Update/ca
      -- 
    ca_1941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_600_inst_ack_1, ack => inputPort_3_Daemon_CP_1763_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	19 
    -- CP-element group 69: 	37 
    -- CP-element group 69: 	43 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_610_Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_610_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_610_sample_start_
      -- 
    rr_1949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(69), ack => EQ_u8_u1_610_inst_req_0); -- 
    inputPort_3_Daemon_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_1763_elements(19) & inputPort_3_Daemon_CP_1763_elements(37) & inputPort_3_Daemon_CP_1763_elements(43);
      gj_inputPort_3_Daemon_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	93 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_610_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_610_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_610_update_start_
      -- 
    cr_1954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(70), ack => EQ_u8_u1_610_inst_req_1); -- 
    inputPort_3_Daemon_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_3_Daemon_CP_1763_elements(93);
      gj_inputPort_3_Daemon_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: marked-successors 
    -- CP-element group 71: 	17 
    -- CP-element group 71: 	33 
    -- CP-element group 71: 	39 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_610_Sample/ra
      -- CP-element group 71: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_610_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_610_sample_completed_
      -- 
    ra_1950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_610_inst_ack_0, ack => inputPort_3_Daemon_CP_1763_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	92 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_610_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_610_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_610_update_completed_
      -- 
    ca_1955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_610_inst_ack_1, ack => inputPort_3_Daemon_CP_1763_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	19 
    -- CP-element group 73: 	37 
    -- CP-element group 73: 	43 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_620_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_620_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_620_Sample/rr
      -- 
    rr_1963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(73), ack => EQ_u8_u1_620_inst_req_0); -- 
    inputPort_3_Daemon_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_1763_elements(19) & inputPort_3_Daemon_CP_1763_elements(37) & inputPort_3_Daemon_CP_1763_elements(43);
      gj_inputPort_3_Daemon_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	99 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_620_Update/cr
      -- CP-element group 74: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_620_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_620_update_start_
      -- 
    cr_1968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(74), ack => EQ_u8_u1_620_inst_req_1); -- 
    inputPort_3_Daemon_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_3_Daemon_CP_1763_elements(99);
      gj_inputPort_3_Daemon_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	17 
    -- CP-element group 75: 	33 
    -- CP-element group 75: 	39 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_620_Sample/ra
      -- CP-element group 75: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_620_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_620_sample_completed_
      -- 
    ra_1964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_620_inst_ack_0, ack => inputPort_3_Daemon_CP_1763_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	98 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_620_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_620_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/EQ_u8_u1_620_Update/ca
      -- 
    ca_1969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_620_inst_ack_1, ack => inputPort_3_Daemon_CP_1763_elements(76)); -- 
    -- CP-element group 77:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	81 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_629_Update/req
      -- CP-element group 77: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_629_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_629_update_start_
      -- 
    req_1982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(77), ack => W_data_to_outport_569_delayed_4_0_627_inst_req_1); -- 
    inputPort_3_Daemon_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_3_Daemon_CP_1763_elements(81);
      gj_inputPort_3_Daemon_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	37 
    -- CP-element group 78: successors 
    -- CP-element group 78: marked-successors 
    -- CP-element group 78: 	33 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_629_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_629_Sample/ack
      -- CP-element group 78: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_629_Sample/$exit
      -- 
    ack_1978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_569_delayed_4_0_627_inst_ack_0, ack => inputPort_3_Daemon_CP_1763_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_629_Update/ack
      -- CP-element group 79: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_629_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_629_update_completed_
      -- 
    ack_1983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_569_delayed_4_0_627_inst_ack_1, ack => inputPort_3_Daemon_CP_1763_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	60 
    -- CP-element group 80: 	79 
    -- CP-element group 80: 	64 
    -- CP-element group 80: marked-predecessors 
    -- CP-element group 80: 	82 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_1_631_Sample/req
      -- CP-element group 80: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_1_631_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_1_631_Sample/$entry
      -- 
    req_1991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(80), ack => WPIPE_noblock_obuf_3_1_631_inst_req_0); -- 
    inputPort_3_Daemon_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_1763_elements(60) & inputPort_3_Daemon_CP_1763_elements(79) & inputPort_3_Daemon_CP_1763_elements(64) & inputPort_3_Daemon_CP_1763_elements(82);
      gj_inputPort_3_Daemon_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81: marked-successors 
    -- CP-element group 81: 	58 
    -- CP-element group 81: 	62 
    -- CP-element group 81: 	77 
    -- CP-element group 81:  members (6) 
      -- CP-element group 81: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_1_631_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_1_631_Sample/ack
      -- CP-element group 81: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_1_631_update_start_
      -- CP-element group 81: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_1_631_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_1_631_Update/req
      -- CP-element group 81: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_1_631_Sample/$exit
      -- 
    ack_1992_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_1_631_inst_ack_0, ack => inputPort_3_Daemon_CP_1763_elements(81)); -- 
    req_1996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(81), ack => WPIPE_noblock_obuf_3_1_631_inst_req_1); -- 
    -- CP-element group 82:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	102 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	80 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_1_631_Update/ack
      -- CP-element group 82: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_1_631_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_1_631_Update/$exit
      -- 
    ack_1997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_1_631_inst_ack_1, ack => inputPort_3_Daemon_CP_1763_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: marked-predecessors 
    -- CP-element group 83: 	87 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_636_update_start_
      -- CP-element group 83: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_636_Update/req
      -- CP-element group 83: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_636_Update/$entry
      -- 
    req_2010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(83), ack => W_data_to_outport_573_delayed_4_0_634_inst_req_1); -- 
    inputPort_3_Daemon_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_3_Daemon_CP_1763_elements(87);
      gj_inputPort_3_Daemon_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	37 
    -- CP-element group 84: successors 
    -- CP-element group 84: marked-successors 
    -- CP-element group 84: 	33 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_636_Sample/ack
      -- CP-element group 84: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_636_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_636_sample_completed_
      -- 
    ack_2006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_573_delayed_4_0_634_inst_ack_0, ack => inputPort_3_Daemon_CP_1763_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_636_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_636_Update/ack
      -- CP-element group 85: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_636_Update/$exit
      -- 
    ack_2011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_573_delayed_4_0_634_inst_ack_1, ack => inputPort_3_Daemon_CP_1763_elements(85)); -- 
    -- CP-element group 86:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: 	68 
    -- CP-element group 86: 	60 
    -- CP-element group 86: marked-predecessors 
    -- CP-element group 86: 	88 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_2_638_Sample/req
      -- CP-element group 86: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_2_638_Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_2_638_sample_start_
      -- 
    req_2019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(86), ack => WPIPE_noblock_obuf_3_2_638_inst_req_0); -- 
    inputPort_3_Daemon_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_1763_elements(85) & inputPort_3_Daemon_CP_1763_elements(68) & inputPort_3_Daemon_CP_1763_elements(60) & inputPort_3_Daemon_CP_1763_elements(88);
      gj_inputPort_3_Daemon_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: marked-successors 
    -- CP-element group 87: 	58 
    -- CP-element group 87: 	66 
    -- CP-element group 87: 	83 
    -- CP-element group 87:  members (6) 
      -- CP-element group 87: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_2_638_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_2_638_Update/req
      -- CP-element group 87: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_2_638_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_2_638_Sample/ack
      -- CP-element group 87: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_2_638_update_start_
      -- CP-element group 87: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_2_638_sample_completed_
      -- 
    ack_2020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_2_638_inst_ack_0, ack => inputPort_3_Daemon_CP_1763_elements(87)); -- 
    req_2024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(87), ack => WPIPE_noblock_obuf_3_2_638_inst_req_1); -- 
    -- CP-element group 88:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	102 
    -- CP-element group 88: marked-successors 
    -- CP-element group 88: 	86 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_2_638_Update/ack
      -- CP-element group 88: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_2_638_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_2_638_update_completed_
      -- 
    ack_2025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_2_638_inst_ack_1, ack => inputPort_3_Daemon_CP_1763_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	93 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_643_update_start_
      -- CP-element group 89: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_643_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_643_Update/req
      -- 
    req_2038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(89), ack => W_data_to_outport_577_delayed_4_0_641_inst_req_1); -- 
    inputPort_3_Daemon_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_3_Daemon_CP_1763_elements(93);
      gj_inputPort_3_Daemon_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	37 
    -- CP-element group 90: successors 
    -- CP-element group 90: marked-successors 
    -- CP-element group 90: 	33 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_643_Sample/ack
      -- CP-element group 90: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_643_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_643_Sample/$exit
      -- 
    ack_2034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_577_delayed_4_0_641_inst_ack_0, ack => inputPort_3_Daemon_CP_1763_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_643_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_643_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_643_Update/ack
      -- 
    ack_2039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_577_delayed_4_0_641_inst_ack_1, ack => inputPort_3_Daemon_CP_1763_elements(91)); -- 
    -- CP-element group 92:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: 	60 
    -- CP-element group 92: 	72 
    -- CP-element group 92: marked-predecessors 
    -- CP-element group 92: 	94 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_3_645_Sample/req
      -- CP-element group 92: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_3_645_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_3_645_sample_start_
      -- 
    req_2047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(92), ack => WPIPE_noblock_obuf_3_3_645_inst_req_0); -- 
    inputPort_3_Daemon_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_1763_elements(91) & inputPort_3_Daemon_CP_1763_elements(60) & inputPort_3_Daemon_CP_1763_elements(72) & inputPort_3_Daemon_CP_1763_elements(94);
      gj_inputPort_3_Daemon_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93: marked-successors 
    -- CP-element group 93: 	58 
    -- CP-element group 93: 	89 
    -- CP-element group 93: 	70 
    -- CP-element group 93:  members (6) 
      -- CP-element group 93: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_3_645_Sample/ack
      -- CP-element group 93: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_3_645_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_3_645_Update/$entry
      -- CP-element group 93: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_3_645_Update/req
      -- CP-element group 93: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_3_645_update_start_
      -- CP-element group 93: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_3_645_sample_completed_
      -- 
    ack_2048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_3_645_inst_ack_0, ack => inputPort_3_Daemon_CP_1763_elements(93)); -- 
    req_2052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(93), ack => WPIPE_noblock_obuf_3_3_645_inst_req_1); -- 
    -- CP-element group 94:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	102 
    -- CP-element group 94: marked-successors 
    -- CP-element group 94: 	92 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_3_645_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_3_645_Update/ack
      -- CP-element group 94: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_3_645_update_completed_
      -- 
    ack_2053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_3_645_inst_ack_1, ack => inputPort_3_Daemon_CP_1763_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: marked-predecessors 
    -- CP-element group 95: 	99 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_650_update_start_
      -- CP-element group 95: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_650_Update/$entry
      -- CP-element group 95: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_650_Update/req
      -- 
    req_2066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(95), ack => W_data_to_outport_581_delayed_4_0_648_inst_req_1); -- 
    inputPort_3_Daemon_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_3_Daemon_CP_1763_elements(99);
      gj_inputPort_3_Daemon_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	37 
    -- CP-element group 96: successors 
    -- CP-element group 96: marked-successors 
    -- CP-element group 96: 	33 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_650_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_650_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_650_Sample/ack
      -- 
    ack_2062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_581_delayed_4_0_648_inst_ack_0, ack => inputPort_3_Daemon_CP_1763_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_650_Update/ack
      -- CP-element group 97: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_650_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/assign_stmt_650_update_completed_
      -- 
    ack_2067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_581_delayed_4_0_648_inst_ack_1, ack => inputPort_3_Daemon_CP_1763_elements(97)); -- 
    -- CP-element group 98:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: 	60 
    -- CP-element group 98: 	76 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	100 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_4_652_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_4_652_Sample/req
      -- CP-element group 98: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_4_652_Sample/$entry
      -- 
    req_2075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(98), ack => WPIPE_noblock_obuf_3_4_652_inst_req_0); -- 
    inputPort_3_Daemon_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_1763_elements(97) & inputPort_3_Daemon_CP_1763_elements(60) & inputPort_3_Daemon_CP_1763_elements(76) & inputPort_3_Daemon_CP_1763_elements(100);
      gj_inputPort_3_Daemon_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: marked-successors 
    -- CP-element group 99: 	58 
    -- CP-element group 99: 	95 
    -- CP-element group 99: 	74 
    -- CP-element group 99:  members (6) 
      -- CP-element group 99: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_4_652_update_start_
      -- CP-element group 99: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_4_652_Sample/ack
      -- CP-element group 99: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_4_652_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_4_652_Update/req
      -- CP-element group 99: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_4_652_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_4_652_Update/$entry
      -- 
    ack_2076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_4_652_inst_ack_0, ack => inputPort_3_Daemon_CP_1763_elements(99)); -- 
    req_2080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_1763_elements(99), ack => WPIPE_noblock_obuf_3_4_652_inst_req_1); -- 
    -- CP-element group 100:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100: marked-successors 
    -- CP-element group 100: 	98 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_4_652_Update/ack
      -- CP-element group 100: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_4_652_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/WPIPE_noblock_obuf_3_4_652_update_completed_
      -- 
    ack_2081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_4_652_inst_ack_1, ack => inputPort_3_Daemon_CP_1763_elements(100)); -- 
    -- CP-element group 101:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	9 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	10 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group inputPort_3_Daemon_CP_1763_elements(101) is a control-delay.
    cp_element_101_delay: control_delay_element  generic map(name => " 101_delay", delay_value => 1)  port map(req => inputPort_3_Daemon_CP_1763_elements(9), ack => inputPort_3_Daemon_CP_1763_elements(101), clk => clk, reset =>reset);
    -- CP-element group 102:  join  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	88 
    -- CP-element group 102: 	100 
    -- CP-element group 102: 	12 
    -- CP-element group 102: 	13 
    -- CP-element group 102: 	94 
    -- CP-element group 102: 	82 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	6 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_518/do_while_stmt_519/do_while_stmt_519_loop_body/$exit
      -- 
    inputPort_3_Daemon_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 39) := "inputPort_3_Daemon_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_1763_elements(88) & inputPort_3_Daemon_CP_1763_elements(100) & inputPort_3_Daemon_CP_1763_elements(12) & inputPort_3_Daemon_CP_1763_elements(13) & inputPort_3_Daemon_CP_1763_elements(94) & inputPort_3_Daemon_CP_1763_elements(82);
      gj_inputPort_3_Daemon_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	5 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_518/do_while_stmt_519/loop_exit/$exit
      -- CP-element group 103: 	 branch_block_stmt_518/do_while_stmt_519/loop_exit/ack
      -- 
    ack_2086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_519_branch_ack_0, ack => inputPort_3_Daemon_CP_1763_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	5 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_518/do_while_stmt_519/loop_taken/ack
      -- CP-element group 104: 	 branch_block_stmt_518/do_while_stmt_519/loop_taken/$exit
      -- 
    ack_2090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_519_branch_ack_1, ack => inputPort_3_Daemon_CP_1763_elements(104)); -- 
    -- CP-element group 105:  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	3 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	1 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_518/do_while_stmt_519/$exit
      -- 
    inputPort_3_Daemon_CP_1763_elements(105) <= inputPort_3_Daemon_CP_1763_elements(3);
    inputPort_3_Daemon_do_while_stmt_519_terminator_2091: loop_terminator -- 
      generic map (name => " inputPort_3_Daemon_do_while_stmt_519_terminator_2091", max_iterations_in_flight =>7) 
      port map(loop_body_exit => inputPort_3_Daemon_CP_1763_elements(6),loop_continue => inputPort_3_Daemon_CP_1763_elements(104),loop_terminate => inputPort_3_Daemon_CP_1763_elements(103),loop_back => inputPort_3_Daemon_CP_1763_elements(4),loop_exit => inputPort_3_Daemon_CP_1763_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_521_phi_seq_1837_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_3_Daemon_CP_1763_elements(22);
      inputPort_3_Daemon_CP_1763_elements(25)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_3_Daemon_CP_1763_elements(25);
      inputPort_3_Daemon_CP_1763_elements(26)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_3_Daemon_CP_1763_elements(27);
      inputPort_3_Daemon_CP_1763_elements(23) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_3_Daemon_CP_1763_elements(20);
      inputPort_3_Daemon_CP_1763_elements(29)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_3_Daemon_CP_1763_elements(31);
      inputPort_3_Daemon_CP_1763_elements(30)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_3_Daemon_CP_1763_elements(32);
      inputPort_3_Daemon_CP_1763_elements(21) <= phi_mux_reqs(1);
      phi_stmt_521_phi_seq_1837 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_521_phi_seq_1837") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_3_Daemon_CP_1763_elements(11), 
          phi_sample_ack => inputPort_3_Daemon_CP_1763_elements(18), 
          phi_update_req => inputPort_3_Daemon_CP_1763_elements(14), 
          phi_update_ack => inputPort_3_Daemon_CP_1763_elements(19), 
          phi_mux_ack => inputPort_3_Daemon_CP_1763_elements(24), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_528_phi_seq_1899_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_3_Daemon_CP_1763_elements(46);
      inputPort_3_Daemon_CP_1763_elements(49)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_3_Daemon_CP_1763_elements(49);
      inputPort_3_Daemon_CP_1763_elements(50)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_3_Daemon_CP_1763_elements(51);
      inputPort_3_Daemon_CP_1763_elements(47) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_3_Daemon_CP_1763_elements(44);
      inputPort_3_Daemon_CP_1763_elements(53)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_3_Daemon_CP_1763_elements(55);
      inputPort_3_Daemon_CP_1763_elements(54)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_3_Daemon_CP_1763_elements(56);
      inputPort_3_Daemon_CP_1763_elements(45) <= phi_mux_reqs(1);
      phi_stmt_528_phi_seq_1899 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_528_phi_seq_1899") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_3_Daemon_CP_1763_elements(40), 
          phi_sample_ack => inputPort_3_Daemon_CP_1763_elements(41), 
          phi_update_req => inputPort_3_Daemon_CP_1763_elements(42), 
          phi_update_ack => inputPort_3_Daemon_CP_1763_elements(43), 
          phi_mux_ack => inputPort_3_Daemon_CP_1763_elements(48), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1788_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= inputPort_3_Daemon_CP_1763_elements(7);
        preds(1)  <= inputPort_3_Daemon_CP_1763_elements(8);
        entry_tmerge_1788 : transition_merge -- 
          generic map(name => " entry_tmerge_1788")
          port map (preds => preds, symbol_out => inputPort_3_Daemon_CP_1763_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal EQ_u8_u1_542_542_delayed_4_0_591 : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_549_549_delayed_4_0_601 : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_556_556_delayed_4_0_611 : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_563_563_delayed_4_0_621 : std_logic_vector(0 downto 0);
    signal RPIPE_in_data_3_527_wire : std_logic_vector(31 downto 0);
    signal R_ONE_1_574_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_16_523_wire_constant : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_561_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_564_wire : std_logic_vector(15 downto 0);
    signal SUB_u8_u8_582_wire : std_logic_vector(7 downto 0);
    signal continue_586 : std_logic_vector(0 downto 0);
    signal count_down_521 : std_logic_vector(15 downto 0);
    signal data_to_outport_569_delayed_4_0_629 : std_logic_vector(32 downto 0);
    signal data_to_outport_573_delayed_4_0_636 : std_logic_vector(32 downto 0);
    signal data_to_outport_577 : std_logic_vector(32 downto 0);
    signal data_to_outport_577_delayed_4_0_643 : std_logic_vector(32 downto 0);
    signal data_to_outport_581_delayed_4_0_650 : std_logic_vector(32 downto 0);
    signal dest_id_543 : std_logic_vector(7 downto 0);
    signal input_word_525 : std_logic_vector(31 downto 0);
    signal konst_530_wire_constant : std_logic_vector(7 downto 0);
    signal konst_537_wire_constant : std_logic_vector(15 downto 0);
    signal konst_560_wire_constant : std_logic_vector(15 downto 0);
    signal konst_563_wire_constant : std_logic_vector(15 downto 0);
    signal konst_579_wire_constant : std_logic_vector(7 downto 0);
    signal konst_581_wire_constant : std_logic_vector(7 downto 0);
    signal konst_589_wire_constant : std_logic_vector(7 downto 0);
    signal konst_599_wire_constant : std_logic_vector(7 downto 0);
    signal konst_609_wire_constant : std_logic_vector(7 downto 0);
    signal konst_619_wire_constant : std_logic_vector(7 downto 0);
    signal konst_666_wire_constant : std_logic_vector(0 downto 0);
    signal last_dest_id_528 : std_logic_vector(7 downto 0);
    signal new_packet_539 : std_logic_vector(0 downto 0);
    signal next_count_down_566 : std_logic_vector(15 downto 0);
    signal next_count_down_566_524_buffered : std_logic_vector(15 downto 0);
    signal next_last_dest_id_572 : std_logic_vector(7 downto 0);
    signal next_last_dest_id_572_531_buffered : std_logic_vector(7 downto 0);
    signal pkt_length_547 : std_logic_vector(15 downto 0);
    signal send_to_1_596 : std_logic_vector(0 downto 0);
    signal send_to_2_606 : std_logic_vector(0 downto 0);
    signal send_to_3_616 : std_logic_vector(0 downto 0);
    signal send_to_4_626 : std_logic_vector(0 downto 0);
    signal seq_id_551 : std_logic_vector(7 downto 0);
    signal type_cast_584_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_ONE_1_574_wire_constant <= "1";
    R_ZERO_16_523_wire_constant <= "0000000000000000";
    konst_530_wire_constant <= "00000000";
    konst_537_wire_constant <= "0000000000000000";
    konst_560_wire_constant <= "0000000000000001";
    konst_563_wire_constant <= "0000000000000001";
    konst_579_wire_constant <= "00000010";
    konst_581_wire_constant <= "00000001";
    konst_589_wire_constant <= "00000001";
    konst_599_wire_constant <= "00000010";
    konst_609_wire_constant <= "00000011";
    konst_619_wire_constant <= "00000100";
    konst_666_wire_constant <= "1";
    type_cast_584_wire_constant <= "1";
    phi_stmt_521: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_16_523_wire_constant & next_count_down_566_524_buffered;
      req <= phi_stmt_521_req_0 & phi_stmt_521_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_521",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_521_ack_0,
          idata => idata,
          odata => count_down_521,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_521
    phi_stmt_528: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= konst_530_wire_constant & next_last_dest_id_572_531_buffered;
      req <= phi_stmt_528_req_0 & phi_stmt_528_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_528",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_528_ack_0,
          idata => idata,
          odata => last_dest_id_528,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_528
    -- flow-through select operator MUX_565_inst
    next_count_down_566 <= SUB_u16_u16_561_wire when (new_packet_539(0) /=  '0') else SUB_u16_u16_564_wire;
    -- flow-through select operator MUX_571_inst
    next_last_dest_id_572 <= dest_id_543 when (new_packet_539(0) /=  '0') else last_dest_id_528;
    -- flow-through slice operator slice_542_inst
    dest_id_543 <= input_word_525(31 downto 24);
    -- flow-through slice operator slice_546_inst
    pkt_length_547 <= input_word_525(23 downto 8);
    -- flow-through slice operator slice_550_inst
    seq_id_551 <= input_word_525(7 downto 0);
    W_data_to_outport_569_delayed_4_0_627_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_data_to_outport_569_delayed_4_0_627_inst_req_0;
      W_data_to_outport_569_delayed_4_0_627_inst_ack_0<= wack(0);
      rreq(0) <= W_data_to_outport_569_delayed_4_0_627_inst_req_1;
      W_data_to_outport_569_delayed_4_0_627_inst_ack_1<= rack(0);
      W_data_to_outport_569_delayed_4_0_627_inst : InterlockBuffer generic map ( -- 
        name => "W_data_to_outport_569_delayed_4_0_627_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 33,
        out_data_width => 33,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => data_to_outport_577,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => data_to_outport_569_delayed_4_0_629,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_data_to_outport_573_delayed_4_0_634_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_data_to_outport_573_delayed_4_0_634_inst_req_0;
      W_data_to_outport_573_delayed_4_0_634_inst_ack_0<= wack(0);
      rreq(0) <= W_data_to_outport_573_delayed_4_0_634_inst_req_1;
      W_data_to_outport_573_delayed_4_0_634_inst_ack_1<= rack(0);
      W_data_to_outport_573_delayed_4_0_634_inst : InterlockBuffer generic map ( -- 
        name => "W_data_to_outport_573_delayed_4_0_634_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 33,
        out_data_width => 33,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => data_to_outport_577,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => data_to_outport_573_delayed_4_0_636,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_data_to_outport_577_delayed_4_0_641_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_data_to_outport_577_delayed_4_0_641_inst_req_0;
      W_data_to_outport_577_delayed_4_0_641_inst_ack_0<= wack(0);
      rreq(0) <= W_data_to_outport_577_delayed_4_0_641_inst_req_1;
      W_data_to_outport_577_delayed_4_0_641_inst_ack_1<= rack(0);
      W_data_to_outport_577_delayed_4_0_641_inst : InterlockBuffer generic map ( -- 
        name => "W_data_to_outport_577_delayed_4_0_641_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 33,
        out_data_width => 33,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => data_to_outport_577,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => data_to_outport_577_delayed_4_0_643,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_data_to_outport_581_delayed_4_0_648_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_data_to_outport_581_delayed_4_0_648_inst_req_0;
      W_data_to_outport_581_delayed_4_0_648_inst_ack_0<= wack(0);
      rreq(0) <= W_data_to_outport_581_delayed_4_0_648_inst_req_1;
      W_data_to_outport_581_delayed_4_0_648_inst_ack_1<= rack(0);
      W_data_to_outport_581_delayed_4_0_648_inst : InterlockBuffer generic map ( -- 
        name => "W_data_to_outport_581_delayed_4_0_648_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 33,
        out_data_width => 33,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => data_to_outport_577,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => data_to_outport_581_delayed_4_0_650,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_count_down_566_524_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_count_down_566_524_buf_req_0;
      next_count_down_566_524_buf_ack_0<= wack(0);
      rreq(0) <= next_count_down_566_524_buf_req_1;
      next_count_down_566_524_buf_ack_1<= rack(0);
      next_count_down_566_524_buf : InterlockBuffer generic map ( -- 
        name => "next_count_down_566_524_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_count_down_566,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_count_down_566_524_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_last_dest_id_572_531_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_last_dest_id_572_531_buf_req_0;
      next_last_dest_id_572_531_buf_ack_0<= wack(0);
      rreq(0) <= next_last_dest_id_572_531_buf_req_1;
      next_last_dest_id_572_531_buf_ack_1<= rack(0);
      next_last_dest_id_572_531_buf : InterlockBuffer generic map ( -- 
        name => "next_last_dest_id_572_531_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_last_dest_id_572,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_last_dest_id_572_531_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_525
    process(RPIPE_in_data_3_527_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := RPIPE_in_data_3_527_wire(31 downto 0);
      input_word_525 <= tmp_var; -- 
    end process;
    do_while_stmt_519_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_666_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_519_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_519_branch_req_0,
          ack0 => do_while_stmt_519_branch_ack_0,
          ack1 => do_while_stmt_519_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- flow through binary operator AND_u1_u1_595_inst
    send_to_1_596 <= (EQ_u8_u1_542_542_delayed_4_0_591 and continue_586);
    -- flow through binary operator AND_u1_u1_605_inst
    send_to_2_606 <= (EQ_u8_u1_549_549_delayed_4_0_601 and continue_586);
    -- flow through binary operator AND_u1_u1_615_inst
    send_to_3_616 <= (EQ_u8_u1_556_556_delayed_4_0_611 and continue_586);
    -- flow through binary operator AND_u1_u1_625_inst
    send_to_4_626 <= (EQ_u8_u1_563_563_delayed_4_0_621 and continue_586);
    -- flow through binary operator CONCAT_u1_u33_576_inst
    process(R_ONE_1_574_wire_constant, input_word_525) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ONE_1_574_wire_constant, input_word_525, tmp_var);
      data_to_outport_577 <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u16_u1_538_inst
    process(count_down_521) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(count_down_521, konst_537_wire_constant, tmp_var);
      new_packet_539 <= tmp_var; --
    end process;
    -- shared split operator group (6) : EQ_u8_u1_590_inst 
    ApIntEq_group_6: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 4);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= next_last_dest_id_572;
      EQ_u8_u1_542_542_delayed_4_0_591 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u8_u1_590_inst_req_0;
      EQ_u8_u1_590_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u8_u1_590_inst_req_1;
      EQ_u8_u1_590_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_6_gI: SplitGuardInterface generic map(name => "ApIntEq_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000001",
          constant_width => 8,
          buffering  => 4,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : EQ_u8_u1_600_inst 
    ApIntEq_group_7: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 4);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= next_last_dest_id_572;
      EQ_u8_u1_549_549_delayed_4_0_601 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u8_u1_600_inst_req_0;
      EQ_u8_u1_600_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u8_u1_600_inst_req_1;
      EQ_u8_u1_600_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_7_gI: SplitGuardInterface generic map(name => "ApIntEq_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000010",
          constant_width => 8,
          buffering  => 4,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : EQ_u8_u1_610_inst 
    ApIntEq_group_8: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 4);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= next_last_dest_id_572;
      EQ_u8_u1_556_556_delayed_4_0_611 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u8_u1_610_inst_req_0;
      EQ_u8_u1_610_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u8_u1_610_inst_req_1;
      EQ_u8_u1_610_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_8_gI: SplitGuardInterface generic map(name => "ApIntEq_group_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_8",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000011",
          constant_width => 8,
          buffering  => 4,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : EQ_u8_u1_620_inst 
    ApIntEq_group_9: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 4);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= next_last_dest_id_572;
      EQ_u8_u1_563_563_delayed_4_0_621 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u8_u1_620_inst_req_0;
      EQ_u8_u1_620_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u8_u1_620_inst_req_1;
      EQ_u8_u1_620_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_9_gI: SplitGuardInterface generic map(name => "ApIntEq_group_9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_9",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000100",
          constant_width => 8,
          buffering  => 4,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- flow through binary operator SUB_u16_u16_561_inst
    SUB_u16_u16_561_wire <= std_logic_vector(unsigned(pkt_length_547) - unsigned(konst_560_wire_constant));
    -- flow through binary operator SUB_u16_u16_564_inst
    SUB_u16_u16_564_wire <= std_logic_vector(unsigned(count_down_521) - unsigned(konst_563_wire_constant));
    -- flow through binary operator SUB_u8_u8_582_inst
    SUB_u8_u8_582_wire <= std_logic_vector(unsigned(next_last_dest_id_572) - unsigned(konst_581_wire_constant));
    -- shared inport operator group (0) : RPIPE_in_data_3_527_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_in_data_3_527_inst_req_0;
      RPIPE_in_data_3_527_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_in_data_3_527_inst_req_1;
      RPIPE_in_data_3_527_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_in_data_3_527_wire <= data_out(31 downto 0);
      in_data_3_read_0_gI: SplitGuardInterface generic map(name => "in_data_3_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      in_data_3_read_0: InputPortRevised -- 
        generic map ( name => "in_data_3_read_0", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => in_data_3_pipe_read_req(0),
          oack => in_data_3_pipe_read_ack(0),
          odata => in_data_3_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_noblock_obuf_3_1_631_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_3_1_631_inst_req_0;
      WPIPE_noblock_obuf_3_1_631_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_3_1_631_inst_req_1;
      WPIPE_noblock_obuf_3_1_631_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_1_596(0);
      data_in <= data_to_outport_569_delayed_4_0_629;
      noblock_obuf_3_1_write_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_1_write_0: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_3_1", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_3_1_pipe_write_req(0),
          oack => noblock_obuf_3_1_pipe_write_ack(0),
          odata => noblock_obuf_3_1_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_noblock_obuf_3_2_638_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_3_2_638_inst_req_0;
      WPIPE_noblock_obuf_3_2_638_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_3_2_638_inst_req_1;
      WPIPE_noblock_obuf_3_2_638_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_2_606(0);
      data_in <= data_to_outport_573_delayed_4_0_636;
      noblock_obuf_3_2_write_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_2_write_1: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_3_2", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_3_2_pipe_write_req(0),
          oack => noblock_obuf_3_2_pipe_write_ack(0),
          odata => noblock_obuf_3_2_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_noblock_obuf_3_3_645_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_3_3_645_inst_req_0;
      WPIPE_noblock_obuf_3_3_645_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_3_3_645_inst_req_1;
      WPIPE_noblock_obuf_3_3_645_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_3_616(0);
      data_in <= data_to_outport_577_delayed_4_0_643;
      noblock_obuf_3_3_write_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_3_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_3_write_2: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_3_3", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_3_3_pipe_write_req(0),
          oack => noblock_obuf_3_3_pipe_write_ack(0),
          odata => noblock_obuf_3_3_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_noblock_obuf_3_4_652_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_3_4_652_inst_req_0;
      WPIPE_noblock_obuf_3_4_652_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_3_4_652_inst_req_1;
      WPIPE_noblock_obuf_3_4_652_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_4_626(0);
      data_in <= data_to_outport_581_delayed_4_0_650;
      noblock_obuf_3_4_write_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_4_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_4_write_3: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_3_4", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_3_4_pipe_write_req(0),
          oack => noblock_obuf_3_4_pipe_write_ack(0),
          odata => noblock_obuf_3_4_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared call operator group (0) : call_updateCounter_expr_585_inst 
    updateCounter_call_group_0: Block -- 
      signal data_in: std_logic_vector(16 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_updateCounter_expr_585_inst_req_0;
      call_updateCounter_expr_585_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_updateCounter_expr_585_inst_req_1;
      call_updateCounter_expr_585_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      updateCounter_call_group_0_gI: SplitGuardInterface generic map(name => "updateCounter_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_579_wire_constant & SUB_u8_u8_582_wire & type_cast_584_wire_constant;
      continue_586 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 17,
        owidth => 17,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => updateCounter_call_reqs(0),
          ackR => updateCounter_call_acks(0),
          dataR => updateCounter_call_data(16 downto 0),
          tagR => updateCounter_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => updateCounter_return_acks(0), -- cross-over
          ackL => updateCounter_return_reqs(0), -- cross-over
          dataL => updateCounter_return_data(0 downto 0),
          tagL => updateCounter_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end inputPort_3_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity inputPort_4_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    in_data_4_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_4_pipe_read_data : in   std_logic_vector(31 downto 0);
    noblock_obuf_4_1_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_1_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_4_2_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_2_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_4_3_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_3_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_4_4_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_4_pipe_write_data : out  std_logic_vector(32 downto 0);
    updateCounter_call_reqs : out  std_logic_vector(0 downto 0);
    updateCounter_call_acks : in   std_logic_vector(0 downto 0);
    updateCounter_call_data : out  std_logic_vector(16 downto 0);
    updateCounter_call_tag  :  out  std_logic_vector(0 downto 0);
    updateCounter_return_reqs : out  std_logic_vector(0 downto 0);
    updateCounter_return_acks : in   std_logic_vector(0 downto 0);
    updateCounter_return_data : in   std_logic_vector(0 downto 0);
    updateCounter_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity inputPort_4_Daemon;
architecture inputPort_4_Daemon_arch of inputPort_4_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal inputPort_4_Daemon_CP_2092_start: Boolean;
  signal inputPort_4_Daemon_CP_2092_symbol: Boolean;
  -- volatile/operator module components. 
  component updateCounter is -- 
    generic (tag_length : integer); 
    port ( -- 
      input_port : in  std_logic_vector(7 downto 0);
      output_port : in  std_logic_vector(7 downto 0);
      up : in  std_logic_vector(0 downto 0);
      continue : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(3 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(1 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(1 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal WPIPE_noblock_obuf_4_2_790_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_4_1_783_inst_req_1 : boolean;
  signal W_data_to_outport_709_delayed_4_0_800_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_4_4_804_inst_req_1 : boolean;
  signal W_data_to_outport_709_delayed_4_0_800_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_4_4_804_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_4_1_783_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_4_3_797_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_4_4_804_inst_ack_0 : boolean;
  signal W_data_to_outport_705_delayed_4_0_793_inst_ack_0 : boolean;
  signal W_data_to_outport_705_delayed_4_0_793_inst_req_0 : boolean;
  signal W_data_to_outport_701_delayed_4_0_786_inst_req_0 : boolean;
  signal W_data_to_outport_701_delayed_4_0_786_inst_ack_0 : boolean;
  signal do_while_stmt_671_branch_ack_0 : boolean;
  signal WPIPE_noblock_obuf_4_2_790_inst_req_1 : boolean;
  signal do_while_stmt_671_branch_ack_1 : boolean;
  signal W_data_to_outport_705_delayed_4_0_793_inst_req_1 : boolean;
  signal W_data_to_outport_701_delayed_4_0_786_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_4_2_790_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_4_3_797_inst_req_1 : boolean;
  signal W_data_to_outport_705_delayed_4_0_793_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_4_3_797_inst_ack_1 : boolean;
  signal W_data_to_outport_709_delayed_4_0_800_inst_req_1 : boolean;
  signal W_data_to_outport_709_delayed_4_0_800_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_4_1_783_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_4_1_783_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_4_3_797_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_4_2_790_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_4_4_804_inst_req_0 : boolean;
  signal W_data_to_outport_701_delayed_4_0_786_inst_ack_1 : boolean;
  signal do_while_stmt_671_branch_req_0 : boolean;
  signal phi_stmt_673_req_1 : boolean;
  signal phi_stmt_673_req_0 : boolean;
  signal phi_stmt_673_ack_0 : boolean;
  signal next_count_down_718_676_buf_req_0 : boolean;
  signal next_count_down_718_676_buf_ack_0 : boolean;
  signal next_count_down_718_676_buf_req_1 : boolean;
  signal next_count_down_718_676_buf_ack_1 : boolean;
  signal RPIPE_in_data_4_679_inst_req_0 : boolean;
  signal RPIPE_in_data_4_679_inst_ack_0 : boolean;
  signal RPIPE_in_data_4_679_inst_req_1 : boolean;
  signal RPIPE_in_data_4_679_inst_ack_1 : boolean;
  signal phi_stmt_680_req_1 : boolean;
  signal phi_stmt_680_req_0 : boolean;
  signal phi_stmt_680_ack_0 : boolean;
  signal next_last_dest_id_724_683_buf_req_0 : boolean;
  signal next_last_dest_id_724_683_buf_ack_0 : boolean;
  signal next_last_dest_id_724_683_buf_req_1 : boolean;
  signal next_last_dest_id_724_683_buf_ack_1 : boolean;
  signal call_updateCounter_expr_737_inst_req_0 : boolean;
  signal call_updateCounter_expr_737_inst_ack_0 : boolean;
  signal call_updateCounter_expr_737_inst_req_1 : boolean;
  signal call_updateCounter_expr_737_inst_ack_1 : boolean;
  signal EQ_u8_u1_742_inst_req_0 : boolean;
  signal EQ_u8_u1_742_inst_ack_0 : boolean;
  signal EQ_u8_u1_742_inst_req_1 : boolean;
  signal EQ_u8_u1_742_inst_ack_1 : boolean;
  signal EQ_u8_u1_752_inst_req_0 : boolean;
  signal EQ_u8_u1_752_inst_ack_0 : boolean;
  signal EQ_u8_u1_752_inst_req_1 : boolean;
  signal EQ_u8_u1_752_inst_ack_1 : boolean;
  signal EQ_u8_u1_762_inst_req_0 : boolean;
  signal EQ_u8_u1_762_inst_ack_0 : boolean;
  signal EQ_u8_u1_762_inst_req_1 : boolean;
  signal EQ_u8_u1_762_inst_ack_1 : boolean;
  signal EQ_u8_u1_772_inst_req_0 : boolean;
  signal EQ_u8_u1_772_inst_ack_0 : boolean;
  signal EQ_u8_u1_772_inst_req_1 : boolean;
  signal EQ_u8_u1_772_inst_ack_1 : boolean;
  signal W_data_to_outport_697_delayed_4_0_779_inst_req_0 : boolean;
  signal W_data_to_outport_697_delayed_4_0_779_inst_ack_0 : boolean;
  signal W_data_to_outport_697_delayed_4_0_779_inst_req_1 : boolean;
  signal W_data_to_outport_697_delayed_4_0_779_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "inputPort_4_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  inputPort_4_Daemon_CP_2092_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "inputPort_4_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_4_Daemon_CP_2092_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= inputPort_4_Daemon_CP_2092_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_4_Daemon_CP_2092_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  inputPort_4_Daemon_CP_2092: Block -- control-path 
    signal inputPort_4_Daemon_CP_2092_elements: BooleanArray(105 downto 0);
    -- 
  begin -- 
    inputPort_4_Daemon_CP_2092_elements(0) <= inputPort_4_Daemon_CP_2092_start;
    inputPort_4_Daemon_CP_2092_symbol <= inputPort_4_Daemon_CP_2092_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_670/$entry
      -- CP-element group 0: 	 branch_block_stmt_670/branch_block_stmt_670__entry__
      -- CP-element group 0: 	 branch_block_stmt_670/do_while_stmt_671__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	105 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_670/$exit
      -- CP-element group 1: 	 branch_block_stmt_670/branch_block_stmt_670__exit__
      -- CP-element group 1: 	 branch_block_stmt_670/do_while_stmt_671__exit__
      -- 
    inputPort_4_Daemon_CP_2092_elements(1) <= inputPort_4_Daemon_CP_2092_elements(105);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_670/do_while_stmt_671/$entry
      -- CP-element group 2: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671__entry__
      -- 
    inputPort_4_Daemon_CP_2092_elements(2) <= inputPort_4_Daemon_CP_2092_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	105 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671__exit__
      -- 
    -- Element group inputPort_4_Daemon_CP_2092_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_670/do_while_stmt_671/loop_back
      -- 
    -- Element group inputPort_4_Daemon_CP_2092_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	103 
    -- CP-element group 5: 	104 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_670/do_while_stmt_671/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_670/do_while_stmt_671/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_670/do_while_stmt_671/condition_done
      -- 
    inputPort_4_Daemon_CP_2092_elements(5) <= inputPort_4_Daemon_CP_2092_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	102 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_670/do_while_stmt_671/loop_body_done
      -- 
    inputPort_4_Daemon_CP_2092_elements(6) <= inputPort_4_Daemon_CP_2092_elements(102);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	20 
    -- CP-element group 7: 	44 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/back_edge_to_loop_body
      -- 
    inputPort_4_Daemon_CP_2092_elements(7) <= inputPort_4_Daemon_CP_2092_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	22 
    -- CP-element group 8: 	46 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/first_time_through_loop_body
      -- 
    inputPort_4_Daemon_CP_2092_elements(8) <= inputPort_4_Daemon_CP_2092_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	17 
    -- CP-element group 9: 	101 
    -- CP-element group 9: 	33 
    -- CP-element group 9: 	38 
    -- CP-element group 9: 	39 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_677_sample_start_
      -- 
    -- Element group inputPort_4_Daemon_CP_2092_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	101 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/condition_evaluated
      -- 
    condition_evaluated_2116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(10), ack => do_while_stmt_671_branch_req_0); -- 
    inputPort_4_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_2092_elements(15) & inputPort_4_Daemon_CP_2092_elements(101);
      gj_inputPort_4_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	16 
    -- CP-element group 11: 	38 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	40 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_673_sample_start__ps
      -- 
    inputPort_4_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_2092_elements(9) & inputPort_4_Daemon_CP_2092_elements(16) & inputPort_4_Daemon_CP_2092_elements(38) & inputPort_4_Daemon_CP_2092_elements(15);
      gj_inputPort_4_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	18 
    -- CP-element group 12: 	36 
    -- CP-element group 12: 	41 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12: 	102 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	16 
    -- CP-element group 12: 	38 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_673_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_677_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_680_sample_completed_
      -- 
    inputPort_4_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_2092_elements(18) & inputPort_4_Daemon_CP_2092_elements(36) & inputPort_4_Daemon_CP_2092_elements(41);
      gj_inputPort_4_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	102 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/aggregated_phi_sample_ack_d
      -- 
    -- Element group inputPort_4_Daemon_CP_2092_elements(13) is a control-delay.
    cp_element_13_delay: control_delay_element  generic map(name => " 13_delay", delay_value => 1)  port map(req => inputPort_4_Daemon_CP_2092_elements(12), ack => inputPort_4_Daemon_CP_2092_elements(13), clk => clk, reset =>reset);
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	17 
    -- CP-element group 14: 	33 
    -- CP-element group 14: 	39 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	35 
    -- CP-element group 14: 	42 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/aggregated_phi_update_req
      -- CP-element group 14: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_673_update_start__ps
      -- 
    inputPort_4_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_2092_elements(17) & inputPort_4_Daemon_CP_2092_elements(33) & inputPort_4_Daemon_CP_2092_elements(39);
      gj_inputPort_4_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	19 
    -- CP-element group 15: 	37 
    -- CP-element group 15: 	43 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/aggregated_phi_update_ack
      -- 
    inputPort_4_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_2092_elements(19) & inputPort_4_Daemon_CP_2092_elements(37) & inputPort_4_Daemon_CP_2092_elements(43);
      gj_inputPort_4_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	11 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_673_sample_start_
      -- 
    inputPort_4_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_2092_elements(9) & inputPort_4_Daemon_CP_2092_elements(12);
      gj_inputPort_4_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	9 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	71 
    -- CP-element group 17: 	67 
    -- CP-element group 17: 	75 
    -- CP-element group 17: 	59 
    -- CP-element group 17: 	63 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	14 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_673_update_start_
      -- 
    inputPort_4_Daemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_2092_elements(9) & inputPort_4_Daemon_CP_2092_elements(71) & inputPort_4_Daemon_CP_2092_elements(67) & inputPort_4_Daemon_CP_2092_elements(75) & inputPort_4_Daemon_CP_2092_elements(59) & inputPort_4_Daemon_CP_2092_elements(63);
      gj_inputPort_4_Daemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_673_sample_completed__ps
      -- 
    -- Element group inputPort_4_Daemon_CP_2092_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: 	65 
    -- CP-element group 19: 	69 
    -- CP-element group 19: 	73 
    -- CP-element group 19: 	57 
    -- CP-element group 19: 	61 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_673_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_673_update_completed__ps
      -- 
    -- Element group inputPort_4_Daemon_CP_2092_elements(19) is bound as output of CP function.
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	7 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_673_loopback_trigger
      -- 
    inputPort_4_Daemon_CP_2092_elements(20) <= inputPort_4_Daemon_CP_2092_elements(7);
    -- CP-element group 21:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_673_loopback_sample_req
      -- CP-element group 21: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_673_loopback_sample_req_ps
      -- 
    phi_stmt_673_loopback_sample_req_2132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_673_loopback_sample_req_2132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(21), ack => phi_stmt_673_req_1); -- 
    -- Element group inputPort_4_Daemon_CP_2092_elements(21) is bound as output of CP function.
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	8 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_673_entry_trigger
      -- 
    inputPort_4_Daemon_CP_2092_elements(22) <= inputPort_4_Daemon_CP_2092_elements(8);
    -- CP-element group 23:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_673_entry_sample_req
      -- CP-element group 23: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_673_entry_sample_req_ps
      -- 
    phi_stmt_673_entry_sample_req_2135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_673_entry_sample_req_2135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(23), ack => phi_stmt_673_req_0); -- 
    -- Element group inputPort_4_Daemon_CP_2092_elements(23) is bound as output of CP function.
    -- CP-element group 24:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_673_phi_mux_ack
      -- CP-element group 24: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_673_phi_mux_ack_ps
      -- 
    phi_stmt_673_phi_mux_ack_2138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_673_ack_0, ack => inputPort_4_Daemon_CP_2092_elements(24)); -- 
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_ZERO_16_675_sample_start__ps
      -- CP-element group 25: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_ZERO_16_675_sample_completed__ps
      -- CP-element group 25: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_ZERO_16_675_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_ZERO_16_675_sample_completed_
      -- 
    -- Element group inputPort_4_Daemon_CP_2092_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_ZERO_16_675_update_start__ps
      -- CP-element group 26: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_ZERO_16_675_update_start_
      -- 
    -- Element group inputPort_4_Daemon_CP_2092_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	28 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_ZERO_16_675_update_completed__ps
      -- 
    inputPort_4_Daemon_CP_2092_elements(27) <= inputPort_4_Daemon_CP_2092_elements(28);
    -- CP-element group 28:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	27 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_ZERO_16_675_update_completed_
      -- 
    -- Element group inputPort_4_Daemon_CP_2092_elements(28) is a control-delay.
    cp_element_28_delay: control_delay_element  generic map(name => " 28_delay", delay_value => 1)  port map(req => inputPort_4_Daemon_CP_2092_elements(26), ack => inputPort_4_Daemon_CP_2092_elements(28), clk => clk, reset =>reset);
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_count_down_676_sample_start__ps
      -- CP-element group 29: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_count_down_676_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_count_down_676_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_count_down_676_Sample/req
      -- 
    req_2159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(29), ack => next_count_down_718_676_buf_req_0); -- 
    -- Element group inputPort_4_Daemon_CP_2092_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_count_down_676_update_start__ps
      -- CP-element group 30: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_count_down_676_update_start_
      -- CP-element group 30: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_count_down_676_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_count_down_676_Update/req
      -- 
    req_2164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(30), ack => next_count_down_718_676_buf_req_1); -- 
    -- Element group inputPort_4_Daemon_CP_2092_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_count_down_676_sample_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_count_down_676_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_count_down_676_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_count_down_676_Sample/ack
      -- 
    ack_2160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_718_676_buf_ack_0, ack => inputPort_4_Daemon_CP_2092_elements(31)); -- 
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_count_down_676_update_completed__ps
      -- CP-element group 32: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_count_down_676_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_count_down_676_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_count_down_676_Update/ack
      -- 
    ack_2165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_718_676_buf_ack_1, ack => inputPort_4_Daemon_CP_2092_elements(32)); -- 
    -- CP-element group 33:  join  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	9 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	78 
    -- CP-element group 33: 	96 
    -- CP-element group 33: 	71 
    -- CP-element group 33: 	84 
    -- CP-element group 33: 	90 
    -- CP-element group 33: 	67 
    -- CP-element group 33: 	75 
    -- CP-element group 33: 	59 
    -- CP-element group 33: 	63 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	14 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_677_update_start_
      -- 
    inputPort_4_Daemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_2092_elements(9) & inputPort_4_Daemon_CP_2092_elements(78) & inputPort_4_Daemon_CP_2092_elements(96) & inputPort_4_Daemon_CP_2092_elements(71) & inputPort_4_Daemon_CP_2092_elements(84) & inputPort_4_Daemon_CP_2092_elements(90) & inputPort_4_Daemon_CP_2092_elements(67) & inputPort_4_Daemon_CP_2092_elements(75) & inputPort_4_Daemon_CP_2092_elements(59) & inputPort_4_Daemon_CP_2092_elements(63);
      gj_inputPort_4_Daemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	11 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	37 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/RPIPE_in_data_4_679_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/RPIPE_in_data_4_679_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/RPIPE_in_data_4_679_Sample/rr
      -- 
    rr_2178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(34), ack => RPIPE_in_data_4_679_inst_req_0); -- 
    inputPort_4_Daemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_2092_elements(11) & inputPort_4_Daemon_CP_2092_elements(37);
      gj_inputPort_4_Daemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	14 
    -- CP-element group 35: 	36 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/RPIPE_in_data_4_679_update_start_
      -- CP-element group 35: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/RPIPE_in_data_4_679_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/RPIPE_in_data_4_679_Update/cr
      -- 
    cr_2183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(35), ack => RPIPE_in_data_4_679_inst_req_1); -- 
    inputPort_4_Daemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_2092_elements(14) & inputPort_4_Daemon_CP_2092_elements(36);
      gj_inputPort_4_Daemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	12 
    -- CP-element group 36: 	35 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/RPIPE_in_data_4_679_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/RPIPE_in_data_4_679_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/RPIPE_in_data_4_679_Sample/ra
      -- 
    ra_2179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_4_679_inst_ack_0, ack => inputPort_4_Daemon_CP_2092_elements(36)); -- 
    -- CP-element group 37:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	15 
    -- CP-element group 37: 	78 
    -- CP-element group 37: 	96 
    -- CP-element group 37: 	84 
    -- CP-element group 37: 	65 
    -- CP-element group 37: 	90 
    -- CP-element group 37: 	69 
    -- CP-element group 37: 	73 
    -- CP-element group 37: 	57 
    -- CP-element group 37: 	61 
    -- CP-element group 37: marked-successors 
    -- CP-element group 37: 	34 
    -- CP-element group 37:  members (16) 
      -- CP-element group 37: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_788_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_802_Sample/req
      -- CP-element group 37: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_802_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_788_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_795_Sample/req
      -- CP-element group 37: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_788_Sample/req
      -- CP-element group 37: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_795_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_802_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_795_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_677_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/RPIPE_in_data_4_679_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/RPIPE_in_data_4_679_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/RPIPE_in_data_4_679_Update/ca
      -- CP-element group 37: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_781_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_781_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_781_Sample/req
      -- 
    ca_2184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_4_679_inst_ack_1, ack => inputPort_4_Daemon_CP_2092_elements(37)); -- 
    req_2362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(37), ack => W_data_to_outport_705_delayed_4_0_793_inst_req_0); -- 
    req_2306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(37), ack => W_data_to_outport_697_delayed_4_0_779_inst_req_0); -- 
    req_2334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(37), ack => W_data_to_outport_701_delayed_4_0_786_inst_req_0); -- 
    req_2390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(37), ack => W_data_to_outport_709_delayed_4_0_800_inst_req_0); -- 
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	9 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	12 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	11 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_680_sample_start_
      -- 
    inputPort_4_Daemon_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_2092_elements(9) & inputPort_4_Daemon_CP_2092_elements(12);
      gj_inputPort_4_Daemon_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  join  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	9 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	71 
    -- CP-element group 39: 	67 
    -- CP-element group 39: 	75 
    -- CP-element group 39: 	59 
    -- CP-element group 39: 	63 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	14 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_680_update_start_
      -- 
    inputPort_4_Daemon_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_2092_elements(9) & inputPort_4_Daemon_CP_2092_elements(71) & inputPort_4_Daemon_CP_2092_elements(67) & inputPort_4_Daemon_CP_2092_elements(75) & inputPort_4_Daemon_CP_2092_elements(59) & inputPort_4_Daemon_CP_2092_elements(63);
      gj_inputPort_4_Daemon_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	11 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_680_sample_start__ps
      -- 
    inputPort_4_Daemon_CP_2092_elements(40) <= inputPort_4_Daemon_CP_2092_elements(11);
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	12 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_680_sample_completed__ps
      -- 
    -- Element group inputPort_4_Daemon_CP_2092_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	14 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_680_update_start__ps
      -- 
    inputPort_4_Daemon_CP_2092_elements(42) <= inputPort_4_Daemon_CP_2092_elements(14);
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	15 
    -- CP-element group 43: 	65 
    -- CP-element group 43: 	69 
    -- CP-element group 43: 	73 
    -- CP-element group 43: 	57 
    -- CP-element group 43: 	61 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_680_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_680_update_completed__ps
      -- 
    -- Element group inputPort_4_Daemon_CP_2092_elements(43) is bound as output of CP function.
    -- CP-element group 44:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	7 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_680_loopback_trigger
      -- 
    inputPort_4_Daemon_CP_2092_elements(44) <= inputPort_4_Daemon_CP_2092_elements(7);
    -- CP-element group 45:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_680_loopback_sample_req
      -- CP-element group 45: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_680_loopback_sample_req_ps
      -- 
    phi_stmt_680_loopback_sample_req_2194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_680_loopback_sample_req_2194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(45), ack => phi_stmt_680_req_1); -- 
    -- Element group inputPort_4_Daemon_CP_2092_elements(45) is bound as output of CP function.
    -- CP-element group 46:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	8 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_680_entry_trigger
      -- 
    inputPort_4_Daemon_CP_2092_elements(46) <= inputPort_4_Daemon_CP_2092_elements(8);
    -- CP-element group 47:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_680_entry_sample_req
      -- CP-element group 47: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_680_entry_sample_req_ps
      -- 
    phi_stmt_680_entry_sample_req_2197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_680_entry_sample_req_2197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(47), ack => phi_stmt_680_req_0); -- 
    -- Element group inputPort_4_Daemon_CP_2092_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_680_phi_mux_ack
      -- CP-element group 48: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/phi_stmt_680_phi_mux_ack_ps
      -- 
    phi_stmt_680_phi_mux_ack_2200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_680_ack_0, ack => inputPort_4_Daemon_CP_2092_elements(48)); -- 
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/konst_682_sample_start__ps
      -- CP-element group 49: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/konst_682_sample_completed__ps
      -- CP-element group 49: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/konst_682_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/konst_682_sample_completed_
      -- 
    -- Element group inputPort_4_Daemon_CP_2092_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (2) 
      -- CP-element group 50: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/konst_682_update_start__ps
      -- CP-element group 50: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/konst_682_update_start_
      -- 
    -- Element group inputPort_4_Daemon_CP_2092_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	52 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/konst_682_update_completed__ps
      -- 
    inputPort_4_Daemon_CP_2092_elements(51) <= inputPort_4_Daemon_CP_2092_elements(52);
    -- CP-element group 52:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	51 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/konst_682_update_completed_
      -- 
    -- Element group inputPort_4_Daemon_CP_2092_elements(52) is a control-delay.
    cp_element_52_delay: control_delay_element  generic map(name => " 52_delay", delay_value => 1)  port map(req => inputPort_4_Daemon_CP_2092_elements(50), ack => inputPort_4_Daemon_CP_2092_elements(52), clk => clk, reset =>reset);
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_last_dest_id_683_sample_start__ps
      -- CP-element group 53: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_last_dest_id_683_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_last_dest_id_683_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_last_dest_id_683_Sample/req
      -- 
    req_2221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(53), ack => next_last_dest_id_724_683_buf_req_0); -- 
    -- Element group inputPort_4_Daemon_CP_2092_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_last_dest_id_683_update_start__ps
      -- CP-element group 54: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_last_dest_id_683_update_start_
      -- CP-element group 54: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_last_dest_id_683_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_last_dest_id_683_Update/req
      -- 
    req_2226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(54), ack => next_last_dest_id_724_683_buf_req_1); -- 
    -- Element group inputPort_4_Daemon_CP_2092_elements(54) is bound as output of CP function.
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_last_dest_id_683_sample_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_last_dest_id_683_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_last_dest_id_683_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_last_dest_id_683_Sample/ack
      -- 
    ack_2222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_724_683_buf_ack_0, ack => inputPort_4_Daemon_CP_2092_elements(55)); -- 
    -- CP-element group 56:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_last_dest_id_683_update_completed__ps
      -- CP-element group 56: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_last_dest_id_683_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_last_dest_id_683_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/R_next_last_dest_id_683_Update/ack
      -- 
    ack_2227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_724_683_buf_ack_1, ack => inputPort_4_Daemon_CP_2092_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	19 
    -- CP-element group 57: 	37 
    -- CP-element group 57: 	43 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/call_updateCounter_expr_737_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/call_updateCounter_expr_737_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/call_updateCounter_expr_737_Sample/req
      -- 
    req_2236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(57), ack => call_updateCounter_expr_737_inst_req_0); -- 
    inputPort_4_Daemon_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_2092_elements(19) & inputPort_4_Daemon_CP_2092_elements(37) & inputPort_4_Daemon_CP_2092_elements(43);
      gj_inputPort_4_Daemon_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	81 
    -- CP-element group 58: 	99 
    -- CP-element group 58: 	87 
    -- CP-element group 58: 	93 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/call_updateCounter_expr_737_update_start_
      -- CP-element group 58: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/call_updateCounter_expr_737_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/call_updateCounter_expr_737_Update/req
      -- 
    req_2241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(58), ack => call_updateCounter_expr_737_inst_req_1); -- 
    inputPort_4_Daemon_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_2092_elements(81) & inputPort_4_Daemon_CP_2092_elements(99) & inputPort_4_Daemon_CP_2092_elements(87) & inputPort_4_Daemon_CP_2092_elements(93);
      gj_inputPort_4_Daemon_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: marked-successors 
    -- CP-element group 59: 	17 
    -- CP-element group 59: 	33 
    -- CP-element group 59: 	39 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/call_updateCounter_expr_737_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/call_updateCounter_expr_737_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/call_updateCounter_expr_737_Sample/ack
      -- 
    ack_2237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_updateCounter_expr_737_inst_ack_0, ack => inputPort_4_Daemon_CP_2092_elements(59)); -- 
    -- CP-element group 60:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	98 
    -- CP-element group 60: 	86 
    -- CP-element group 60: 	92 
    -- CP-element group 60: 	80 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/call_updateCounter_expr_737_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/call_updateCounter_expr_737_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/call_updateCounter_expr_737_Update/ack
      -- 
    ack_2242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_updateCounter_expr_737_inst_ack_1, ack => inputPort_4_Daemon_CP_2092_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	19 
    -- CP-element group 61: 	37 
    -- CP-element group 61: 	43 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_742_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_742_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_742_Sample/rr
      -- 
    rr_2250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(61), ack => EQ_u8_u1_742_inst_req_0); -- 
    inputPort_4_Daemon_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_2092_elements(19) & inputPort_4_Daemon_CP_2092_elements(37) & inputPort_4_Daemon_CP_2092_elements(43);
      gj_inputPort_4_Daemon_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	81 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_742_update_start_
      -- CP-element group 62: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_742_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_742_Update/cr
      -- 
    cr_2255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(62), ack => EQ_u8_u1_742_inst_req_1); -- 
    inputPort_4_Daemon_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_4_Daemon_CP_2092_elements(81);
      gj_inputPort_4_Daemon_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	17 
    -- CP-element group 63: 	33 
    -- CP-element group 63: 	39 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_742_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_742_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_742_Sample/ra
      -- 
    ra_2251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_742_inst_ack_0, ack => inputPort_4_Daemon_CP_2092_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	80 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_742_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_742_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_742_Update/ca
      -- 
    ca_2256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_742_inst_ack_1, ack => inputPort_4_Daemon_CP_2092_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	19 
    -- CP-element group 65: 	37 
    -- CP-element group 65: 	43 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_752_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_752_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_752_Sample/rr
      -- 
    rr_2264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(65), ack => EQ_u8_u1_752_inst_req_0); -- 
    inputPort_4_Daemon_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_2092_elements(19) & inputPort_4_Daemon_CP_2092_elements(37) & inputPort_4_Daemon_CP_2092_elements(43);
      gj_inputPort_4_Daemon_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	87 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_752_update_start_
      -- CP-element group 66: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_752_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_752_Update/cr
      -- 
    cr_2269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(66), ack => EQ_u8_u1_752_inst_req_1); -- 
    inputPort_4_Daemon_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_4_Daemon_CP_2092_elements(87);
      gj_inputPort_4_Daemon_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	17 
    -- CP-element group 67: 	33 
    -- CP-element group 67: 	39 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_752_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_752_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_752_Sample/ra
      -- 
    ra_2265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_752_inst_ack_0, ack => inputPort_4_Daemon_CP_2092_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	86 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_752_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_752_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_752_Update/ca
      -- 
    ca_2270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_752_inst_ack_1, ack => inputPort_4_Daemon_CP_2092_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	19 
    -- CP-element group 69: 	37 
    -- CP-element group 69: 	43 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_762_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_762_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_762_Sample/rr
      -- 
    rr_2278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(69), ack => EQ_u8_u1_762_inst_req_0); -- 
    inputPort_4_Daemon_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_2092_elements(19) & inputPort_4_Daemon_CP_2092_elements(37) & inputPort_4_Daemon_CP_2092_elements(43);
      gj_inputPort_4_Daemon_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	93 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_762_update_start_
      -- CP-element group 70: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_762_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_762_Update/cr
      -- 
    cr_2283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(70), ack => EQ_u8_u1_762_inst_req_1); -- 
    inputPort_4_Daemon_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_4_Daemon_CP_2092_elements(93);
      gj_inputPort_4_Daemon_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: marked-successors 
    -- CP-element group 71: 	17 
    -- CP-element group 71: 	33 
    -- CP-element group 71: 	39 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_762_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_762_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_762_Sample/ra
      -- 
    ra_2279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_762_inst_ack_0, ack => inputPort_4_Daemon_CP_2092_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	92 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_762_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_762_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_762_Update/ca
      -- 
    ca_2284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_762_inst_ack_1, ack => inputPort_4_Daemon_CP_2092_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	19 
    -- CP-element group 73: 	37 
    -- CP-element group 73: 	43 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_772_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_772_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_772_Sample/rr
      -- 
    rr_2292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(73), ack => EQ_u8_u1_772_inst_req_0); -- 
    inputPort_4_Daemon_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_2092_elements(19) & inputPort_4_Daemon_CP_2092_elements(37) & inputPort_4_Daemon_CP_2092_elements(43);
      gj_inputPort_4_Daemon_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	99 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_772_update_start_
      -- CP-element group 74: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_772_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_772_Update/cr
      -- 
    cr_2297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(74), ack => EQ_u8_u1_772_inst_req_1); -- 
    inputPort_4_Daemon_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_4_Daemon_CP_2092_elements(99);
      gj_inputPort_4_Daemon_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	17 
    -- CP-element group 75: 	33 
    -- CP-element group 75: 	39 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_772_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_772_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_772_Sample/ra
      -- 
    ra_2293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_772_inst_ack_0, ack => inputPort_4_Daemon_CP_2092_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	98 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_772_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_772_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/EQ_u8_u1_772_Update/ca
      -- 
    ca_2298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_772_inst_ack_1, ack => inputPort_4_Daemon_CP_2092_elements(76)); -- 
    -- CP-element group 77:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	81 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_781_update_start_
      -- CP-element group 77: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_781_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_781_Update/req
      -- 
    req_2311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(77), ack => W_data_to_outport_697_delayed_4_0_779_inst_req_1); -- 
    inputPort_4_Daemon_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_4_Daemon_CP_2092_elements(81);
      gj_inputPort_4_Daemon_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	37 
    -- CP-element group 78: successors 
    -- CP-element group 78: marked-successors 
    -- CP-element group 78: 	33 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_781_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_781_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_781_Sample/ack
      -- 
    ack_2307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_697_delayed_4_0_779_inst_ack_0, ack => inputPort_4_Daemon_CP_2092_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_781_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_781_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_781_Update/ack
      -- 
    ack_2312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_697_delayed_4_0_779_inst_ack_1, ack => inputPort_4_Daemon_CP_2092_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	64 
    -- CP-element group 80: 	79 
    -- CP-element group 80: 	60 
    -- CP-element group 80: marked-predecessors 
    -- CP-element group 80: 	82 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_1_783_Sample/req
      -- CP-element group 80: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_1_783_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_1_783_sample_start_
      -- 
    req_2320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(80), ack => WPIPE_noblock_obuf_4_1_783_inst_req_0); -- 
    inputPort_4_Daemon_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_2092_elements(64) & inputPort_4_Daemon_CP_2092_elements(79) & inputPort_4_Daemon_CP_2092_elements(60) & inputPort_4_Daemon_CP_2092_elements(82);
      gj_inputPort_4_Daemon_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81: marked-successors 
    -- CP-element group 81: 	77 
    -- CP-element group 81: 	58 
    -- CP-element group 81: 	62 
    -- CP-element group 81:  members (6) 
      -- CP-element group 81: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_1_783_Update/req
      -- CP-element group 81: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_1_783_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_1_783_Sample/ack
      -- CP-element group 81: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_1_783_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_1_783_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_1_783_update_start_
      -- 
    ack_2321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_1_783_inst_ack_0, ack => inputPort_4_Daemon_CP_2092_elements(81)); -- 
    req_2325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(81), ack => WPIPE_noblock_obuf_4_1_783_inst_req_1); -- 
    -- CP-element group 82:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	102 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	80 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_1_783_Update/ack
      -- CP-element group 82: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_1_783_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_1_783_update_completed_
      -- 
    ack_2326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_1_783_inst_ack_1, ack => inputPort_4_Daemon_CP_2092_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: marked-predecessors 
    -- CP-element group 83: 	87 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_788_update_start_
      -- CP-element group 83: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_788_Update/$entry
      -- CP-element group 83: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_788_Update/req
      -- 
    req_2339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(83), ack => W_data_to_outport_701_delayed_4_0_786_inst_req_1); -- 
    inputPort_4_Daemon_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_4_Daemon_CP_2092_elements(87);
      gj_inputPort_4_Daemon_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	37 
    -- CP-element group 84: successors 
    -- CP-element group 84: marked-successors 
    -- CP-element group 84: 	33 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_788_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_788_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_788_Sample/ack
      -- 
    ack_2335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_701_delayed_4_0_786_inst_ack_0, ack => inputPort_4_Daemon_CP_2092_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_788_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_788_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_788_Update/ack
      -- 
    ack_2340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_701_delayed_4_0_786_inst_ack_1, ack => inputPort_4_Daemon_CP_2092_elements(85)); -- 
    -- CP-element group 86:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: 	68 
    -- CP-element group 86: 	60 
    -- CP-element group 86: marked-predecessors 
    -- CP-element group 86: 	88 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_2_790_Sample/req
      -- CP-element group 86: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_2_790_Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_2_790_sample_start_
      -- 
    req_2348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(86), ack => WPIPE_noblock_obuf_4_2_790_inst_req_0); -- 
    inputPort_4_Daemon_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_2092_elements(85) & inputPort_4_Daemon_CP_2092_elements(68) & inputPort_4_Daemon_CP_2092_elements(60) & inputPort_4_Daemon_CP_2092_elements(88);
      gj_inputPort_4_Daemon_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: marked-successors 
    -- CP-element group 87: 	83 
    -- CP-element group 87: 	66 
    -- CP-element group 87: 	58 
    -- CP-element group 87:  members (6) 
      -- CP-element group 87: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_2_790_Sample/ack
      -- CP-element group 87: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_2_790_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_2_790_Update/req
      -- CP-element group 87: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_2_790_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_2_790_update_start_
      -- CP-element group 87: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_2_790_sample_completed_
      -- 
    ack_2349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_2_790_inst_ack_0, ack => inputPort_4_Daemon_CP_2092_elements(87)); -- 
    req_2353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(87), ack => WPIPE_noblock_obuf_4_2_790_inst_req_1); -- 
    -- CP-element group 88:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	102 
    -- CP-element group 88: marked-successors 
    -- CP-element group 88: 	86 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_2_790_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_2_790_Update/ack
      -- CP-element group 88: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_2_790_update_completed_
      -- 
    ack_2354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_2_790_inst_ack_1, ack => inputPort_4_Daemon_CP_2092_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	93 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_795_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_795_Update/req
      -- CP-element group 89: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_795_update_start_
      -- 
    req_2367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(89), ack => W_data_to_outport_705_delayed_4_0_793_inst_req_1); -- 
    inputPort_4_Daemon_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_4_Daemon_CP_2092_elements(93);
      gj_inputPort_4_Daemon_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	37 
    -- CP-element group 90: successors 
    -- CP-element group 90: marked-successors 
    -- CP-element group 90: 	33 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_795_Sample/ack
      -- CP-element group 90: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_795_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_795_sample_completed_
      -- 
    ack_2363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_705_delayed_4_0_793_inst_ack_0, ack => inputPort_4_Daemon_CP_2092_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_795_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_795_Update/ack
      -- CP-element group 91: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_795_update_completed_
      -- 
    ack_2368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_705_delayed_4_0_793_inst_ack_1, ack => inputPort_4_Daemon_CP_2092_elements(91)); -- 
    -- CP-element group 92:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	72 
    -- CP-element group 92: 	91 
    -- CP-element group 92: 	60 
    -- CP-element group 92: marked-predecessors 
    -- CP-element group 92: 	94 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_3_797_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_3_797_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_3_797_Sample/req
      -- 
    req_2376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(92), ack => WPIPE_noblock_obuf_4_3_797_inst_req_0); -- 
    inputPort_4_Daemon_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_2092_elements(72) & inputPort_4_Daemon_CP_2092_elements(91) & inputPort_4_Daemon_CP_2092_elements(60) & inputPort_4_Daemon_CP_2092_elements(94);
      gj_inputPort_4_Daemon_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93: marked-successors 
    -- CP-element group 93: 	70 
    -- CP-element group 93: 	89 
    -- CP-element group 93: 	58 
    -- CP-element group 93:  members (6) 
      -- CP-element group 93: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_3_797_Update/$entry
      -- CP-element group 93: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_3_797_Sample/ack
      -- CP-element group 93: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_3_797_Update/req
      -- CP-element group 93: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_3_797_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_3_797_update_start_
      -- CP-element group 93: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_3_797_Sample/$exit
      -- 
    ack_2377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_3_797_inst_ack_0, ack => inputPort_4_Daemon_CP_2092_elements(93)); -- 
    req_2381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(93), ack => WPIPE_noblock_obuf_4_3_797_inst_req_1); -- 
    -- CP-element group 94:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	102 
    -- CP-element group 94: marked-successors 
    -- CP-element group 94: 	92 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_3_797_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_3_797_Update/ack
      -- CP-element group 94: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_3_797_update_completed_
      -- 
    ack_2382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_3_797_inst_ack_1, ack => inputPort_4_Daemon_CP_2092_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: marked-predecessors 
    -- CP-element group 95: 	99 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_802_Update/$entry
      -- CP-element group 95: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_802_Update/req
      -- CP-element group 95: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_802_update_start_
      -- 
    req_2395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(95), ack => W_data_to_outport_709_delayed_4_0_800_inst_req_1); -- 
    inputPort_4_Daemon_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= inputPort_4_Daemon_CP_2092_elements(99);
      gj_inputPort_4_Daemon_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	37 
    -- CP-element group 96: successors 
    -- CP-element group 96: marked-successors 
    -- CP-element group 96: 	33 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_802_Sample/ack
      -- CP-element group 96: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_802_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_802_sample_completed_
      -- 
    ack_2391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_709_delayed_4_0_800_inst_ack_0, ack => inputPort_4_Daemon_CP_2092_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_802_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_802_Update/ack
      -- CP-element group 97: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/assign_stmt_802_update_completed_
      -- 
    ack_2396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_to_outport_709_delayed_4_0_800_inst_ack_1, ack => inputPort_4_Daemon_CP_2092_elements(97)); -- 
    -- CP-element group 98:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: 	76 
    -- CP-element group 98: 	60 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	100 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_4_804_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_4_804_Sample/req
      -- CP-element group 98: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_4_804_Sample/$entry
      -- 
    req_2404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(98), ack => WPIPE_noblock_obuf_4_4_804_inst_req_0); -- 
    inputPort_4_Daemon_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_2092_elements(97) & inputPort_4_Daemon_CP_2092_elements(76) & inputPort_4_Daemon_CP_2092_elements(60) & inputPort_4_Daemon_CP_2092_elements(100);
      gj_inputPort_4_Daemon_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: marked-successors 
    -- CP-element group 99: 	74 
    -- CP-element group 99: 	95 
    -- CP-element group 99: 	58 
    -- CP-element group 99:  members (6) 
      -- CP-element group 99: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_4_804_Update/req
      -- CP-element group 99: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_4_804_Sample/ack
      -- CP-element group 99: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_4_804_Update/$entry
      -- CP-element group 99: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_4_804_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_4_804_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_4_804_update_start_
      -- 
    ack_2405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_4_804_inst_ack_0, ack => inputPort_4_Daemon_CP_2092_elements(99)); -- 
    req_2409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_2092_elements(99), ack => WPIPE_noblock_obuf_4_4_804_inst_req_1); -- 
    -- CP-element group 100:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100: marked-successors 
    -- CP-element group 100: 	98 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_4_804_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_4_804_Update/ack
      -- CP-element group 100: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/WPIPE_noblock_obuf_4_4_804_update_completed_
      -- 
    ack_2410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_4_804_inst_ack_1, ack => inputPort_4_Daemon_CP_2092_elements(100)); -- 
    -- CP-element group 101:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	9 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	10 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group inputPort_4_Daemon_CP_2092_elements(101) is a control-delay.
    cp_element_101_delay: control_delay_element  generic map(name => " 101_delay", delay_value => 1)  port map(req => inputPort_4_Daemon_CP_2092_elements(9), ack => inputPort_4_Daemon_CP_2092_elements(101), clk => clk, reset =>reset);
    -- CP-element group 102:  join  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	12 
    -- CP-element group 102: 	13 
    -- CP-element group 102: 	100 
    -- CP-element group 102: 	88 
    -- CP-element group 102: 	82 
    -- CP-element group 102: 	94 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	6 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_670/do_while_stmt_671/do_while_stmt_671_loop_body/$exit
      -- 
    inputPort_4_Daemon_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 39) := "inputPort_4_Daemon_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_2092_elements(12) & inputPort_4_Daemon_CP_2092_elements(13) & inputPort_4_Daemon_CP_2092_elements(100) & inputPort_4_Daemon_CP_2092_elements(88) & inputPort_4_Daemon_CP_2092_elements(82) & inputPort_4_Daemon_CP_2092_elements(94);
      gj_inputPort_4_Daemon_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	5 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_670/do_while_stmt_671/loop_exit/$exit
      -- CP-element group 103: 	 branch_block_stmt_670/do_while_stmt_671/loop_exit/ack
      -- 
    ack_2415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_671_branch_ack_0, ack => inputPort_4_Daemon_CP_2092_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	5 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_670/do_while_stmt_671/loop_taken/$exit
      -- CP-element group 104: 	 branch_block_stmt_670/do_while_stmt_671/loop_taken/ack
      -- 
    ack_2419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_671_branch_ack_1, ack => inputPort_4_Daemon_CP_2092_elements(104)); -- 
    -- CP-element group 105:  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	3 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	1 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_670/do_while_stmt_671/$exit
      -- 
    inputPort_4_Daemon_CP_2092_elements(105) <= inputPort_4_Daemon_CP_2092_elements(3);
    inputPort_4_Daemon_do_while_stmt_671_terminator_2420: loop_terminator -- 
      generic map (name => " inputPort_4_Daemon_do_while_stmt_671_terminator_2420", max_iterations_in_flight =>7) 
      port map(loop_body_exit => inputPort_4_Daemon_CP_2092_elements(6),loop_continue => inputPort_4_Daemon_CP_2092_elements(104),loop_terminate => inputPort_4_Daemon_CP_2092_elements(103),loop_back => inputPort_4_Daemon_CP_2092_elements(4),loop_exit => inputPort_4_Daemon_CP_2092_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_673_phi_seq_2166_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_4_Daemon_CP_2092_elements(22);
      inputPort_4_Daemon_CP_2092_elements(25)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_4_Daemon_CP_2092_elements(25);
      inputPort_4_Daemon_CP_2092_elements(26)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_4_Daemon_CP_2092_elements(27);
      inputPort_4_Daemon_CP_2092_elements(23) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_4_Daemon_CP_2092_elements(20);
      inputPort_4_Daemon_CP_2092_elements(29)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_4_Daemon_CP_2092_elements(31);
      inputPort_4_Daemon_CP_2092_elements(30)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_4_Daemon_CP_2092_elements(32);
      inputPort_4_Daemon_CP_2092_elements(21) <= phi_mux_reqs(1);
      phi_stmt_673_phi_seq_2166 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_673_phi_seq_2166") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_4_Daemon_CP_2092_elements(11), 
          phi_sample_ack => inputPort_4_Daemon_CP_2092_elements(18), 
          phi_update_req => inputPort_4_Daemon_CP_2092_elements(14), 
          phi_update_ack => inputPort_4_Daemon_CP_2092_elements(19), 
          phi_mux_ack => inputPort_4_Daemon_CP_2092_elements(24), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_680_phi_seq_2228_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_4_Daemon_CP_2092_elements(46);
      inputPort_4_Daemon_CP_2092_elements(49)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_4_Daemon_CP_2092_elements(49);
      inputPort_4_Daemon_CP_2092_elements(50)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_4_Daemon_CP_2092_elements(51);
      inputPort_4_Daemon_CP_2092_elements(47) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_4_Daemon_CP_2092_elements(44);
      inputPort_4_Daemon_CP_2092_elements(53)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_4_Daemon_CP_2092_elements(55);
      inputPort_4_Daemon_CP_2092_elements(54)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_4_Daemon_CP_2092_elements(56);
      inputPort_4_Daemon_CP_2092_elements(45) <= phi_mux_reqs(1);
      phi_stmt_680_phi_seq_2228 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_680_phi_seq_2228") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_4_Daemon_CP_2092_elements(40), 
          phi_sample_ack => inputPort_4_Daemon_CP_2092_elements(41), 
          phi_update_req => inputPort_4_Daemon_CP_2092_elements(42), 
          phi_update_ack => inputPort_4_Daemon_CP_2092_elements(43), 
          phi_mux_ack => inputPort_4_Daemon_CP_2092_elements(48), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_2117_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= inputPort_4_Daemon_CP_2092_elements(7);
        preds(1)  <= inputPort_4_Daemon_CP_2092_elements(8);
        entry_tmerge_2117 : transition_merge -- 
          generic map(name => " entry_tmerge_2117")
          port map (preds => preds, symbol_out => inputPort_4_Daemon_CP_2092_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal EQ_u8_u1_670_670_delayed_4_0_743 : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_677_677_delayed_4_0_753 : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_684_684_delayed_4_0_763 : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_691_691_delayed_4_0_773 : std_logic_vector(0 downto 0);
    signal RPIPE_in_data_4_679_wire : std_logic_vector(31 downto 0);
    signal R_ONE_1_726_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_16_675_wire_constant : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_713_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_716_wire : std_logic_vector(15 downto 0);
    signal SUB_u8_u8_734_wire : std_logic_vector(7 downto 0);
    signal continue_738 : std_logic_vector(0 downto 0);
    signal count_down_673 : std_logic_vector(15 downto 0);
    signal data_to_outport_697_delayed_4_0_781 : std_logic_vector(32 downto 0);
    signal data_to_outport_701_delayed_4_0_788 : std_logic_vector(32 downto 0);
    signal data_to_outport_705_delayed_4_0_795 : std_logic_vector(32 downto 0);
    signal data_to_outport_709_delayed_4_0_802 : std_logic_vector(32 downto 0);
    signal data_to_outport_729 : std_logic_vector(32 downto 0);
    signal dest_id_695 : std_logic_vector(7 downto 0);
    signal input_word_677 : std_logic_vector(31 downto 0);
    signal konst_682_wire_constant : std_logic_vector(7 downto 0);
    signal konst_689_wire_constant : std_logic_vector(15 downto 0);
    signal konst_712_wire_constant : std_logic_vector(15 downto 0);
    signal konst_715_wire_constant : std_logic_vector(15 downto 0);
    signal konst_731_wire_constant : std_logic_vector(7 downto 0);
    signal konst_733_wire_constant : std_logic_vector(7 downto 0);
    signal konst_741_wire_constant : std_logic_vector(7 downto 0);
    signal konst_751_wire_constant : std_logic_vector(7 downto 0);
    signal konst_761_wire_constant : std_logic_vector(7 downto 0);
    signal konst_771_wire_constant : std_logic_vector(7 downto 0);
    signal konst_818_wire_constant : std_logic_vector(0 downto 0);
    signal last_dest_id_680 : std_logic_vector(7 downto 0);
    signal new_packet_691 : std_logic_vector(0 downto 0);
    signal next_count_down_718 : std_logic_vector(15 downto 0);
    signal next_count_down_718_676_buffered : std_logic_vector(15 downto 0);
    signal next_last_dest_id_724 : std_logic_vector(7 downto 0);
    signal next_last_dest_id_724_683_buffered : std_logic_vector(7 downto 0);
    signal pkt_length_699 : std_logic_vector(15 downto 0);
    signal send_to_1_748 : std_logic_vector(0 downto 0);
    signal send_to_2_758 : std_logic_vector(0 downto 0);
    signal send_to_3_768 : std_logic_vector(0 downto 0);
    signal send_to_4_778 : std_logic_vector(0 downto 0);
    signal seq_id_703 : std_logic_vector(7 downto 0);
    signal type_cast_736_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_ONE_1_726_wire_constant <= "1";
    R_ZERO_16_675_wire_constant <= "0000000000000000";
    konst_682_wire_constant <= "00000000";
    konst_689_wire_constant <= "0000000000000000";
    konst_712_wire_constant <= "0000000000000001";
    konst_715_wire_constant <= "0000000000000001";
    konst_731_wire_constant <= "00000011";
    konst_733_wire_constant <= "00000001";
    konst_741_wire_constant <= "00000001";
    konst_751_wire_constant <= "00000010";
    konst_761_wire_constant <= "00000011";
    konst_771_wire_constant <= "00000100";
    konst_818_wire_constant <= "1";
    type_cast_736_wire_constant <= "1";
    phi_stmt_673: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_16_675_wire_constant & next_count_down_718_676_buffered;
      req <= phi_stmt_673_req_0 & phi_stmt_673_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_673",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_673_ack_0,
          idata => idata,
          odata => count_down_673,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_673
    phi_stmt_680: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= konst_682_wire_constant & next_last_dest_id_724_683_buffered;
      req <= phi_stmt_680_req_0 & phi_stmt_680_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_680",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_680_ack_0,
          idata => idata,
          odata => last_dest_id_680,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_680
    -- flow-through select operator MUX_717_inst
    next_count_down_718 <= SUB_u16_u16_713_wire when (new_packet_691(0) /=  '0') else SUB_u16_u16_716_wire;
    -- flow-through select operator MUX_723_inst
    next_last_dest_id_724 <= dest_id_695 when (new_packet_691(0) /=  '0') else last_dest_id_680;
    -- flow-through slice operator slice_694_inst
    dest_id_695 <= input_word_677(31 downto 24);
    -- flow-through slice operator slice_698_inst
    pkt_length_699 <= input_word_677(23 downto 8);
    -- flow-through slice operator slice_702_inst
    seq_id_703 <= input_word_677(7 downto 0);
    W_data_to_outport_697_delayed_4_0_779_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_data_to_outport_697_delayed_4_0_779_inst_req_0;
      W_data_to_outport_697_delayed_4_0_779_inst_ack_0<= wack(0);
      rreq(0) <= W_data_to_outport_697_delayed_4_0_779_inst_req_1;
      W_data_to_outport_697_delayed_4_0_779_inst_ack_1<= rack(0);
      W_data_to_outport_697_delayed_4_0_779_inst : InterlockBuffer generic map ( -- 
        name => "W_data_to_outport_697_delayed_4_0_779_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 33,
        out_data_width => 33,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => data_to_outport_729,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => data_to_outport_697_delayed_4_0_781,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_data_to_outport_701_delayed_4_0_786_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_data_to_outport_701_delayed_4_0_786_inst_req_0;
      W_data_to_outport_701_delayed_4_0_786_inst_ack_0<= wack(0);
      rreq(0) <= W_data_to_outport_701_delayed_4_0_786_inst_req_1;
      W_data_to_outport_701_delayed_4_0_786_inst_ack_1<= rack(0);
      W_data_to_outport_701_delayed_4_0_786_inst : InterlockBuffer generic map ( -- 
        name => "W_data_to_outport_701_delayed_4_0_786_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 33,
        out_data_width => 33,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => data_to_outport_729,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => data_to_outport_701_delayed_4_0_788,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_data_to_outport_705_delayed_4_0_793_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_data_to_outport_705_delayed_4_0_793_inst_req_0;
      W_data_to_outport_705_delayed_4_0_793_inst_ack_0<= wack(0);
      rreq(0) <= W_data_to_outport_705_delayed_4_0_793_inst_req_1;
      W_data_to_outport_705_delayed_4_0_793_inst_ack_1<= rack(0);
      W_data_to_outport_705_delayed_4_0_793_inst : InterlockBuffer generic map ( -- 
        name => "W_data_to_outport_705_delayed_4_0_793_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 33,
        out_data_width => 33,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => data_to_outport_729,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => data_to_outport_705_delayed_4_0_795,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_data_to_outport_709_delayed_4_0_800_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_data_to_outport_709_delayed_4_0_800_inst_req_0;
      W_data_to_outport_709_delayed_4_0_800_inst_ack_0<= wack(0);
      rreq(0) <= W_data_to_outport_709_delayed_4_0_800_inst_req_1;
      W_data_to_outport_709_delayed_4_0_800_inst_ack_1<= rack(0);
      W_data_to_outport_709_delayed_4_0_800_inst : InterlockBuffer generic map ( -- 
        name => "W_data_to_outport_709_delayed_4_0_800_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 33,
        out_data_width => 33,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => data_to_outport_729,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => data_to_outport_709_delayed_4_0_802,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_count_down_718_676_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_count_down_718_676_buf_req_0;
      next_count_down_718_676_buf_ack_0<= wack(0);
      rreq(0) <= next_count_down_718_676_buf_req_1;
      next_count_down_718_676_buf_ack_1<= rack(0);
      next_count_down_718_676_buf : InterlockBuffer generic map ( -- 
        name => "next_count_down_718_676_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_count_down_718,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_count_down_718_676_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_last_dest_id_724_683_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_last_dest_id_724_683_buf_req_0;
      next_last_dest_id_724_683_buf_ack_0<= wack(0);
      rreq(0) <= next_last_dest_id_724_683_buf_req_1;
      next_last_dest_id_724_683_buf_ack_1<= rack(0);
      next_last_dest_id_724_683_buf : InterlockBuffer generic map ( -- 
        name => "next_last_dest_id_724_683_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_last_dest_id_724,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_last_dest_id_724_683_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_677
    process(RPIPE_in_data_4_679_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := RPIPE_in_data_4_679_wire(31 downto 0);
      input_word_677 <= tmp_var; -- 
    end process;
    do_while_stmt_671_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_818_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_671_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_671_branch_req_0,
          ack0 => do_while_stmt_671_branch_ack_0,
          ack1 => do_while_stmt_671_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- flow through binary operator AND_u1_u1_747_inst
    send_to_1_748 <= (EQ_u8_u1_670_670_delayed_4_0_743 and continue_738);
    -- flow through binary operator AND_u1_u1_757_inst
    send_to_2_758 <= (EQ_u8_u1_677_677_delayed_4_0_753 and continue_738);
    -- flow through binary operator AND_u1_u1_767_inst
    send_to_3_768 <= (EQ_u8_u1_684_684_delayed_4_0_763 and continue_738);
    -- flow through binary operator AND_u1_u1_777_inst
    send_to_4_778 <= (EQ_u8_u1_691_691_delayed_4_0_773 and continue_738);
    -- flow through binary operator CONCAT_u1_u33_728_inst
    process(R_ONE_1_726_wire_constant, input_word_677) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ONE_1_726_wire_constant, input_word_677, tmp_var);
      data_to_outport_729 <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u16_u1_690_inst
    process(count_down_673) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(count_down_673, konst_689_wire_constant, tmp_var);
      new_packet_691 <= tmp_var; --
    end process;
    -- shared split operator group (6) : EQ_u8_u1_742_inst 
    ApIntEq_group_6: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 4);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= next_last_dest_id_724;
      EQ_u8_u1_670_670_delayed_4_0_743 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u8_u1_742_inst_req_0;
      EQ_u8_u1_742_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u8_u1_742_inst_req_1;
      EQ_u8_u1_742_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_6_gI: SplitGuardInterface generic map(name => "ApIntEq_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000001",
          constant_width => 8,
          buffering  => 4,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : EQ_u8_u1_752_inst 
    ApIntEq_group_7: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 4);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= next_last_dest_id_724;
      EQ_u8_u1_677_677_delayed_4_0_753 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u8_u1_752_inst_req_0;
      EQ_u8_u1_752_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u8_u1_752_inst_req_1;
      EQ_u8_u1_752_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_7_gI: SplitGuardInterface generic map(name => "ApIntEq_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000010",
          constant_width => 8,
          buffering  => 4,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : EQ_u8_u1_762_inst 
    ApIntEq_group_8: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 4);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= next_last_dest_id_724;
      EQ_u8_u1_684_684_delayed_4_0_763 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u8_u1_762_inst_req_0;
      EQ_u8_u1_762_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u8_u1_762_inst_req_1;
      EQ_u8_u1_762_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_8_gI: SplitGuardInterface generic map(name => "ApIntEq_group_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_8",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000011",
          constant_width => 8,
          buffering  => 4,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : EQ_u8_u1_772_inst 
    ApIntEq_group_9: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 4);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= next_last_dest_id_724;
      EQ_u8_u1_691_691_delayed_4_0_773 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u8_u1_772_inst_req_0;
      EQ_u8_u1_772_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u8_u1_772_inst_req_1;
      EQ_u8_u1_772_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_9_gI: SplitGuardInterface generic map(name => "ApIntEq_group_9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_9",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000100",
          constant_width => 8,
          buffering  => 4,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- flow through binary operator SUB_u16_u16_713_inst
    SUB_u16_u16_713_wire <= std_logic_vector(unsigned(pkt_length_699) - unsigned(konst_712_wire_constant));
    -- flow through binary operator SUB_u16_u16_716_inst
    SUB_u16_u16_716_wire <= std_logic_vector(unsigned(count_down_673) - unsigned(konst_715_wire_constant));
    -- flow through binary operator SUB_u8_u8_734_inst
    SUB_u8_u8_734_wire <= std_logic_vector(unsigned(next_last_dest_id_724) - unsigned(konst_733_wire_constant));
    -- shared inport operator group (0) : RPIPE_in_data_4_679_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_in_data_4_679_inst_req_0;
      RPIPE_in_data_4_679_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_in_data_4_679_inst_req_1;
      RPIPE_in_data_4_679_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_in_data_4_679_wire <= data_out(31 downto 0);
      in_data_4_read_0_gI: SplitGuardInterface generic map(name => "in_data_4_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      in_data_4_read_0: InputPortRevised -- 
        generic map ( name => "in_data_4_read_0", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => in_data_4_pipe_read_req(0),
          oack => in_data_4_pipe_read_ack(0),
          odata => in_data_4_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_noblock_obuf_4_1_783_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_4_1_783_inst_req_0;
      WPIPE_noblock_obuf_4_1_783_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_4_1_783_inst_req_1;
      WPIPE_noblock_obuf_4_1_783_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_1_748(0);
      data_in <= data_to_outport_697_delayed_4_0_781;
      noblock_obuf_4_1_write_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_1_write_0: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_4_1", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_4_1_pipe_write_req(0),
          oack => noblock_obuf_4_1_pipe_write_ack(0),
          odata => noblock_obuf_4_1_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_noblock_obuf_4_2_790_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_4_2_790_inst_req_0;
      WPIPE_noblock_obuf_4_2_790_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_4_2_790_inst_req_1;
      WPIPE_noblock_obuf_4_2_790_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_2_758(0);
      data_in <= data_to_outport_701_delayed_4_0_788;
      noblock_obuf_4_2_write_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_2_write_1: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_4_2", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_4_2_pipe_write_req(0),
          oack => noblock_obuf_4_2_pipe_write_ack(0),
          odata => noblock_obuf_4_2_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_noblock_obuf_4_3_797_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_4_3_797_inst_req_0;
      WPIPE_noblock_obuf_4_3_797_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_4_3_797_inst_req_1;
      WPIPE_noblock_obuf_4_3_797_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_3_768(0);
      data_in <= data_to_outport_705_delayed_4_0_795;
      noblock_obuf_4_3_write_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_3_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_3_write_2: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_4_3", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_4_3_pipe_write_req(0),
          oack => noblock_obuf_4_3_pipe_write_ack(0),
          odata => noblock_obuf_4_3_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_noblock_obuf_4_4_804_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_4_4_804_inst_req_0;
      WPIPE_noblock_obuf_4_4_804_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_4_4_804_inst_req_1;
      WPIPE_noblock_obuf_4_4_804_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_4_778(0);
      data_in <= data_to_outport_709_delayed_4_0_802;
      noblock_obuf_4_4_write_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_4_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_4_write_3: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_4_4", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_4_4_pipe_write_req(0),
          oack => noblock_obuf_4_4_pipe_write_ack(0),
          odata => noblock_obuf_4_4_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared call operator group (0) : call_updateCounter_expr_737_inst 
    updateCounter_call_group_0: Block -- 
      signal data_in: std_logic_vector(16 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_updateCounter_expr_737_inst_req_0;
      call_updateCounter_expr_737_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_updateCounter_expr_737_inst_req_1;
      call_updateCounter_expr_737_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      updateCounter_call_group_0_gI: SplitGuardInterface generic map(name => "updateCounter_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_731_wire_constant & SUB_u8_u8_734_wire & type_cast_736_wire_constant;
      continue_738 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 17,
        owidth => 17,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => updateCounter_call_reqs(0),
          ackR => updateCounter_call_acks(0),
          dataR => updateCounter_call_data(16 downto 0),
          tagR => updateCounter_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => updateCounter_return_acks(0), -- cross-over
          ackL => updateCounter_return_reqs(0), -- cross-over
          dataL => updateCounter_return_data(0 downto 0),
          tagL => updateCounter_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end inputPort_4_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity outputPort_1_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    noblock_obuf_4_1_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_1_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_2_1_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_1_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_1_1_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_1_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_3_1_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_1_pipe_read_data : in   std_logic_vector(32 downto 0);
    out_data_1_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_data_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_data_1_pipe_write_data : out  std_logic_vector(31 downto 0);
    updateCounter_call_reqs : out  std_logic_vector(0 downto 0);
    updateCounter_call_acks : in   std_logic_vector(0 downto 0);
    updateCounter_call_data : out  std_logic_vector(16 downto 0);
    updateCounter_call_tag  :  out  std_logic_vector(0 downto 0);
    updateCounter_return_reqs : out  std_logic_vector(0 downto 0);
    updateCounter_return_acks : in   std_logic_vector(0 downto 0);
    updateCounter_return_data : in   std_logic_vector(0 downto 0);
    updateCounter_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity outputPort_1_Daemon;
architecture outputPort_1_Daemon_arch of outputPort_1_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal outputPort_1_Daemon_CP_2424_start: Boolean;
  signal outputPort_1_Daemon_CP_2424_symbol: Boolean;
  -- volatile/operator module components. 
  component updateCounter is -- 
    generic (tag_length : integer); 
    port ( -- 
      input_port : in  std_logic_vector(7 downto 0);
      output_port : in  std_logic_vector(7 downto 0);
      up : in  std_logic_vector(0 downto 0);
      continue : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(3 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(1 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(1 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component prioritySelect_Volatile is -- 
    port ( -- 
      down_counter : in  std_logic_vector(7 downto 0);
      active_packet : in  std_logic_vector(2 downto 0);
      priority_index : in  std_logic_vector(1 downto 0);
      p1_valid : in  std_logic_vector(0 downto 0);
      p2_valid : in  std_logic_vector(0 downto 0);
      p3_valid : in  std_logic_vector(0 downto 0);
      p4_valid : in  std_logic_vector(0 downto 0);
      next_active_packet : out  std_logic_vector(2 downto 0);
      next_priority_index : out  std_logic_vector(1 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal RPIPE_noblock_obuf_1_1_1053_inst_req_0 : boolean;
  signal phi_stmt_1059_ack_0 : boolean;
  signal RPIPE_noblock_obuf_1_1_1053_inst_ack_1 : boolean;
  signal RPIPE_noblock_obuf_2_1_1058_inst_ack_1 : boolean;
  signal phi_stmt_1059_req_0 : boolean;
  signal RPIPE_noblock_obuf_1_1_1053_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_3_1_1063_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_3_1_1063_inst_req_0 : boolean;
  signal phi_stmt_1054_req_1 : boolean;
  signal phi_stmt_1054_req_0 : boolean;
  signal RPIPE_noblock_obuf_3_1_1063_inst_ack_1 : boolean;
  signal RPIPE_noblock_obuf_2_1_1058_inst_req_0 : boolean;
  signal phi_stmt_1054_ack_0 : boolean;
  signal phi_stmt_1059_req_1 : boolean;
  signal RPIPE_noblock_obuf_2_1_1058_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_2_1_1058_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_3_1_1063_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_1_1_1053_inst_req_1 : boolean;
  signal do_while_stmt_1043_branch_req_0 : boolean;
  signal phi_stmt_1045_req_1 : boolean;
  signal phi_stmt_1045_req_0 : boolean;
  signal phi_stmt_1045_ack_0 : boolean;
  signal next_down_counter_1237_1048_buf_req_0 : boolean;
  signal next_down_counter_1237_1048_buf_ack_0 : boolean;
  signal next_down_counter_1237_1048_buf_req_1 : boolean;
  signal next_down_counter_1237_1048_buf_ack_1 : boolean;
  signal phi_stmt_1049_req_1 : boolean;
  signal phi_stmt_1049_req_0 : boolean;
  signal phi_stmt_1049_ack_0 : boolean;
  signal phi_stmt_1064_req_1 : boolean;
  signal phi_stmt_1064_req_0 : boolean;
  signal phi_stmt_1064_ack_0 : boolean;
  signal RPIPE_noblock_obuf_4_1_1068_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_4_1_1068_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_4_1_1068_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_4_1_1068_inst_ack_1 : boolean;
  signal phi_stmt_1069_req_1 : boolean;
  signal phi_stmt_1069_req_0 : boolean;
  signal phi_stmt_1069_ack_0 : boolean;
  signal next_active_packet_1179_1072_buf_req_0 : boolean;
  signal next_active_packet_1179_1072_buf_ack_0 : boolean;
  signal next_active_packet_1179_1072_buf_req_1 : boolean;
  signal next_active_packet_1179_1072_buf_ack_1 : boolean;
  signal phi_stmt_1073_req_1 : boolean;
  signal phi_stmt_1073_req_0 : boolean;
  signal phi_stmt_1073_ack_0 : boolean;
  signal next_active_packet_length_1224_1076_buf_req_0 : boolean;
  signal next_active_packet_length_1224_1076_buf_ack_0 : boolean;
  signal next_active_packet_length_1224_1076_buf_req_1 : boolean;
  signal next_active_packet_length_1224_1076_buf_ack_1 : boolean;
  signal phi_stmt_1077_req_1 : boolean;
  signal phi_stmt_1077_req_0 : boolean;
  signal phi_stmt_1077_ack_0 : boolean;
  signal next_priority_index_1179_1080_buf_req_0 : boolean;
  signal next_priority_index_1179_1080_buf_ack_0 : boolean;
  signal next_priority_index_1179_1080_buf_req_1 : boolean;
  signal next_priority_index_1179_1080_buf_ack_1 : boolean;
  signal call_stmt_1108_call_req_0 : boolean;
  signal call_stmt_1108_call_ack_0 : boolean;
  signal call_stmt_1108_call_req_1 : boolean;
  signal call_stmt_1108_call_ack_1 : boolean;
  signal WPIPE_out_data_1_1333_inst_req_0 : boolean;
  signal WPIPE_out_data_1_1333_inst_ack_0 : boolean;
  signal WPIPE_out_data_1_1333_inst_req_1 : boolean;
  signal WPIPE_out_data_1_1333_inst_ack_1 : boolean;
  signal do_while_stmt_1043_branch_ack_0 : boolean;
  signal do_while_stmt_1043_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "outputPort_1_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  outputPort_1_Daemon_CP_2424_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "outputPort_1_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_1_Daemon_CP_2424_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= outputPort_1_Daemon_CP_2424_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_1_Daemon_CP_2424_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  outputPort_1_Daemon_CP_2424: Block -- control-path 
    signal outputPort_1_Daemon_CP_2424_elements: BooleanArray(185 downto 0);
    -- 
  begin -- 
    outputPort_1_Daemon_CP_2424_elements(0) <= outputPort_1_Daemon_CP_2424_start;
    outputPort_1_Daemon_CP_2424_symbol <= outputPort_1_Daemon_CP_2424_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1042/$entry
      -- CP-element group 0: 	 branch_block_stmt_1042/branch_block_stmt_1042__entry__
      -- CP-element group 0: 	 branch_block_stmt_1042/do_while_stmt_1043__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	185 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1042/$exit
      -- CP-element group 1: 	 branch_block_stmt_1042/branch_block_stmt_1042__exit__
      -- CP-element group 1: 	 branch_block_stmt_1042/do_while_stmt_1043__exit__
      -- 
    outputPort_1_Daemon_CP_2424_elements(1) <= outputPort_1_Daemon_CP_2424_elements(185);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1042/do_while_stmt_1043/$entry
      -- CP-element group 2: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043__entry__
      -- 
    outputPort_1_Daemon_CP_2424_elements(2) <= outputPort_1_Daemon_CP_2424_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	185 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043__exit__
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1042/do_while_stmt_1043/loop_back
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	183 
    -- CP-element group 5: 	184 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1042/do_while_stmt_1043/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1042/do_while_stmt_1043/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1042/do_while_stmt_1043/loop_taken/$entry
      -- 
    outputPort_1_Daemon_CP_2424_elements(5) <= outputPort_1_Daemon_CP_2424_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	182 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1042/do_while_stmt_1043/loop_body_done
      -- 
    outputPort_1_Daemon_CP_2424_elements(6) <= outputPort_1_Daemon_CP_2424_elements(182);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	142 
    -- CP-element group 7: 	123 
    -- CP-element group 7: 	161 
    -- CP-element group 7: 	22 
    -- CP-element group 7: 	41 
    -- CP-element group 7: 	104 
    -- CP-element group 7: 	62 
    -- CP-element group 7: 	83 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/back_edge_to_loop_body
      -- 
    outputPort_1_Daemon_CP_2424_elements(7) <= outputPort_1_Daemon_CP_2424_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	106 
    -- CP-element group 8: 	144 
    -- CP-element group 8: 	125 
    -- CP-element group 8: 	163 
    -- CP-element group 8: 	24 
    -- CP-element group 8: 	43 
    -- CP-element group 8: 	64 
    -- CP-element group 8: 	85 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/first_time_through_loop_body
      -- 
    outputPort_1_Daemon_CP_2424_elements(8) <= outputPort_1_Daemon_CP_2424_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	181 
    -- CP-element group 9: 	136 
    -- CP-element group 9: 	99 
    -- CP-element group 9: 	98 
    -- CP-element group 9: 	137 
    -- CP-element group 9: 	119 
    -- CP-element group 9: 	120 
    -- CP-element group 9: 	155 
    -- CP-element group 9: 	156 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	17 
    -- CP-element group 9: 	35 
    -- CP-element group 9: 	36 
    -- CP-element group 9: 	56 
    -- CP-element group 9: 	57 
    -- CP-element group 9: 	77 
    -- CP-element group 9: 	78 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/loop_body_start
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	181 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/condition_evaluated
      -- 
    condition_evaluated_2448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(10), ack => do_while_stmt_1043_branch_req_0); -- 
    outputPort_1_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(181) & outputPort_1_Daemon_CP_2424_elements(15);
      gj_outputPort_1_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	136 
    -- CP-element group 11: 	98 
    -- CP-element group 11: 	119 
    -- CP-element group 11: 	155 
    -- CP-element group 11: 	16 
    -- CP-element group 11: 	35 
    -- CP-element group 11: 	56 
    -- CP-element group 11: 	77 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	157 
    -- CP-element group 11: 	138 
    -- CP-element group 11: 	100 
    -- CP-element group 11: 	18 
    -- CP-element group 11: 	37 
    -- CP-element group 11: 	58 
    -- CP-element group 11: 	79 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1069_sample_start__ps
      -- 
    outputPort_1_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 1);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(136) & outputPort_1_Daemon_CP_2424_elements(98) & outputPort_1_Daemon_CP_2424_elements(119) & outputPort_1_Daemon_CP_2424_elements(155) & outputPort_1_Daemon_CP_2424_elements(16) & outputPort_1_Daemon_CP_2424_elements(35) & outputPort_1_Daemon_CP_2424_elements(56) & outputPort_1_Daemon_CP_2424_elements(77) & outputPort_1_Daemon_CP_2424_elements(15);
      gj_outputPort_1_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	121 
    -- CP-element group 12: 	158 
    -- CP-element group 12: 	139 
    -- CP-element group 12: 	101 
    -- CP-element group 12: 	19 
    -- CP-element group 12: 	38 
    -- CP-element group 12: 	59 
    -- CP-element group 12: 	80 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	182 
    -- CP-element group 12: 	13 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	136 
    -- CP-element group 12: 	98 
    -- CP-element group 12: 	119 
    -- CP-element group 12: 	155 
    -- CP-element group 12: 	16 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	56 
    -- CP-element group 12: 	77 
    -- CP-element group 12:  members (9) 
      -- CP-element group 12: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1059_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1054_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1064_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1045_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1049_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1069_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1073_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1077_sample_completed_
      -- 
    outputPort_1_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(121) & outputPort_1_Daemon_CP_2424_elements(158) & outputPort_1_Daemon_CP_2424_elements(139) & outputPort_1_Daemon_CP_2424_elements(101) & outputPort_1_Daemon_CP_2424_elements(19) & outputPort_1_Daemon_CP_2424_elements(38) & outputPort_1_Daemon_CP_2424_elements(59) & outputPort_1_Daemon_CP_2424_elements(80);
      gj_outputPort_1_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	182 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/aggregated_phi_sample_ack_d
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(13) is a control-delay.
    cp_element_13_delay: control_delay_element  generic map(name => " 13_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_2424_elements(12), ack => outputPort_1_Daemon_CP_2424_elements(13), clk => clk, reset =>reset);
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	99 
    -- CP-element group 14: 	137 
    -- CP-element group 14: 	120 
    -- CP-element group 14: 	156 
    -- CP-element group 14: 	17 
    -- CP-element group 14: 	36 
    -- CP-element group 14: 	57 
    -- CP-element group 14: 	78 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	159 
    -- CP-element group 14: 	140 
    -- CP-element group 14: 	102 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	39 
    -- CP-element group 14: 	60 
    -- CP-element group 14: 	81 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/aggregated_phi_update_req
      -- CP-element group 14: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1069_update_start__ps
      -- 
    outputPort_1_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(99) & outputPort_1_Daemon_CP_2424_elements(137) & outputPort_1_Daemon_CP_2424_elements(120) & outputPort_1_Daemon_CP_2424_elements(156) & outputPort_1_Daemon_CP_2424_elements(17) & outputPort_1_Daemon_CP_2424_elements(36) & outputPort_1_Daemon_CP_2424_elements(57) & outputPort_1_Daemon_CP_2424_elements(78);
      gj_outputPort_1_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	122 
    -- CP-element group 15: 	141 
    -- CP-element group 15: 	160 
    -- CP-element group 15: 	21 
    -- CP-element group 15: 	40 
    -- CP-element group 15: 	103 
    -- CP-element group 15: 	61 
    -- CP-element group 15: 	82 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/aggregated_phi_update_ack
      -- 
    outputPort_1_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 7);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(122) & outputPort_1_Daemon_CP_2424_elements(141) & outputPort_1_Daemon_CP_2424_elements(160) & outputPort_1_Daemon_CP_2424_elements(21) & outputPort_1_Daemon_CP_2424_elements(40) & outputPort_1_Daemon_CP_2424_elements(103) & outputPort_1_Daemon_CP_2424_elements(61) & outputPort_1_Daemon_CP_2424_elements(82);
      gj_outputPort_1_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	11 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1045_sample_start_
      -- 
    outputPort_1_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(9) & outputPort_1_Daemon_CP_2424_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	9 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	176 
    -- CP-element group 17: 	179 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	14 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1045_update_start_
      -- 
    outputPort_1_Daemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(9) & outputPort_1_Daemon_CP_2424_elements(176) & outputPort_1_Daemon_CP_2424_elements(179);
      gj_outputPort_1_Daemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	11 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1045_sample_start__ps
      -- 
    outputPort_1_Daemon_CP_2424_elements(18) <= outputPort_1_Daemon_CP_2424_elements(11);
    -- CP-element group 19:  join  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	12 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1045_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(19) is bound as output of CP function.
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	14 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1045_update_start__ps
      -- 
    outputPort_1_Daemon_CP_2424_elements(20) <= outputPort_1_Daemon_CP_2424_elements(14);
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	178 
    -- CP-element group 21: 	174 
    -- CP-element group 21: 	15 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1045_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1045_update_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(21) is bound as output of CP function.
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	7 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1045_loopback_trigger
      -- 
    outputPort_1_Daemon_CP_2424_elements(22) <= outputPort_1_Daemon_CP_2424_elements(7);
    -- CP-element group 23:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1045_loopback_sample_req
      -- CP-element group 23: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1045_loopback_sample_req_ps
      -- 
    phi_stmt_1045_loopback_sample_req_2464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1045_loopback_sample_req_2464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(23), ack => phi_stmt_1045_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(23) is bound as output of CP function.
    -- CP-element group 24:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	8 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1045_entry_trigger
      -- 
    outputPort_1_Daemon_CP_2424_elements(24) <= outputPort_1_Daemon_CP_2424_elements(8);
    -- CP-element group 25:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1045_entry_sample_req
      -- CP-element group 25: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1045_entry_sample_req_ps
      -- 
    phi_stmt_1045_entry_sample_req_2467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1045_entry_sample_req_2467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(25), ack => phi_stmt_1045_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1045_phi_mux_ack
      -- CP-element group 26: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1045_phi_mux_ack_ps
      -- 
    phi_stmt_1045_phi_mux_ack_2470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1045_ack_0, ack => outputPort_1_Daemon_CP_2424_elements(26)); -- 
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_8_1047_sample_start__ps
      -- CP-element group 27: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_8_1047_sample_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_8_1047_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_8_1047_sample_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_8_1047_update_start__ps
      -- CP-element group 28: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_8_1047_update_start_
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	30 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_8_1047_update_completed__ps
      -- 
    outputPort_1_Daemon_CP_2424_elements(29) <= outputPort_1_Daemon_CP_2424_elements(30);
    -- CP-element group 30:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	29 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_8_1047_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(30) is a control-delay.
    cp_element_30_delay: control_delay_element  generic map(name => " 30_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_2424_elements(28), ack => outputPort_1_Daemon_CP_2424_elements(30), clk => clk, reset =>reset);
    -- CP-element group 31:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_down_counter_1048_sample_start__ps
      -- CP-element group 31: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_down_counter_1048_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_down_counter_1048_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_down_counter_1048_Sample/req
      -- 
    req_2491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(31), ack => next_down_counter_1237_1048_buf_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_down_counter_1048_update_start__ps
      -- CP-element group 32: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_down_counter_1048_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_down_counter_1048_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_down_counter_1048_Update/req
      -- 
    req_2496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(32), ack => next_down_counter_1237_1048_buf_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_down_counter_1048_sample_completed__ps
      -- CP-element group 33: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_down_counter_1048_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_down_counter_1048_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_down_counter_1048_Sample/ack
      -- 
    ack_2492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_1237_1048_buf_ack_0, ack => outputPort_1_Daemon_CP_2424_elements(33)); -- 
    -- CP-element group 34:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_down_counter_1048_update_completed__ps
      -- CP-element group 34: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_down_counter_1048_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_down_counter_1048_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_down_counter_1048_Update/ack
      -- 
    ack_2497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_1237_1048_buf_ack_1, ack => outputPort_1_Daemon_CP_2424_elements(34)); -- 
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	12 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	11 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1049_sample_start_
      -- 
    outputPort_1_Daemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(9) & outputPort_1_Daemon_CP_2424_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	9 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	176 
    -- CP-element group 36: 	179 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	14 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1049_update_start_
      -- 
    outputPort_1_Daemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(9) & outputPort_1_Daemon_CP_2424_elements(176) & outputPort_1_Daemon_CP_2424_elements(179);
      gj_outputPort_1_Daemon_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	11 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1049_sample_start__ps
      -- 
    outputPort_1_Daemon_CP_2424_elements(37) <= outputPort_1_Daemon_CP_2424_elements(11);
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	12 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1049_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(38) is bound as output of CP function.
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	14 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1049_update_start__ps
      -- 
    outputPort_1_Daemon_CP_2424_elements(39) <= outputPort_1_Daemon_CP_2424_elements(14);
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	178 
    -- CP-element group 40: 	174 
    -- CP-element group 40: 	15 
    -- CP-element group 40:  members (2) 
      -- CP-element group 40: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1049_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1049_update_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(40) is bound as output of CP function.
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	7 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1049_loopback_trigger
      -- 
    outputPort_1_Daemon_CP_2424_elements(41) <= outputPort_1_Daemon_CP_2424_elements(7);
    -- CP-element group 42:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1049_loopback_sample_req
      -- CP-element group 42: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1049_loopback_sample_req_ps
      -- 
    phi_stmt_1049_loopback_sample_req_2508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1049_loopback_sample_req_2508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(42), ack => phi_stmt_1049_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(42) is bound as output of CP function.
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	8 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1049_entry_trigger
      -- 
    outputPort_1_Daemon_CP_2424_elements(43) <= outputPort_1_Daemon_CP_2424_elements(8);
    -- CP-element group 44:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1049_entry_sample_req
      -- CP-element group 44: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1049_entry_sample_req_ps
      -- 
    phi_stmt_1049_entry_sample_req_2511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1049_entry_sample_req_2511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(44), ack => phi_stmt_1049_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(44) is bound as output of CP function.
    -- CP-element group 45:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1049_phi_mux_ack
      -- CP-element group 45: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1049_phi_mux_ack_ps
      -- 
    phi_stmt_1049_phi_mux_ack_2514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1049_ack_0, ack => outputPort_1_Daemon_CP_2424_elements(45)); -- 
    -- CP-element group 46:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (4) 
      -- CP-element group 46: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1051_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1051_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1051_sample_start__ps
      -- CP-element group 46: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1051_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1051_update_start_
      -- CP-element group 47: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1051_update_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	49 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1051_update_completed__ps
      -- 
    outputPort_1_Daemon_CP_2424_elements(48) <= outputPort_1_Daemon_CP_2424_elements(49);
    -- CP-element group 49:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	48 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1051_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(49) is a control-delay.
    cp_element_49_delay: control_delay_element  generic map(name => " 49_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_2424_elements(47), ack => outputPort_1_Daemon_CP_2424_elements(49), clk => clk, reset =>reset);
    -- CP-element group 50:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_1_1_1053_sample_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_1_1_1053_update_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(51) is bound as output of CP function.
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	55 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_1_1_1053_Sample/rr
      -- CP-element group 52: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_1_1_1053_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_1_1_1053_Sample/$entry
      -- 
    rr_2535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(52), ack => RPIPE_noblock_obuf_1_1_1053_inst_req_0); -- 
    outputPort_1_Daemon_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(50) & outputPort_1_Daemon_CP_2424_elements(55);
      gj_outputPort_1_Daemon_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: 	54 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_1_1_1053_update_start_
      -- CP-element group 53: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_1_1_1053_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_1_1_1053_Update/cr
      -- 
    cr_2540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(53), ack => RPIPE_noblock_obuf_1_1_1053_inst_req_1); -- 
    outputPort_1_Daemon_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(51) & outputPort_1_Daemon_CP_2424_elements(54);
      gj_outputPort_1_Daemon_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	53 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_1_1_1053_sample_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_1_1_1053_Sample/ra
      -- CP-element group 54: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_1_1_1053_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_1_1_1053_Sample/$exit
      -- 
    ra_2536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_1_1053_inst_ack_0, ack => outputPort_1_Daemon_CP_2424_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: marked-successors 
    -- CP-element group 55: 	52 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_1_1_1053_Update/ca
      -- CP-element group 55: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_1_1_1053_update_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_1_1_1053_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_1_1_1053_update_completed_
      -- 
    ca_2541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_1_1053_inst_ack_1, ack => outputPort_1_Daemon_CP_2424_elements(55)); -- 
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	9 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	12 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	11 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1054_sample_start_
      -- 
    outputPort_1_Daemon_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(9) & outputPort_1_Daemon_CP_2424_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  join  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	9 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	176 
    -- CP-element group 57: 	179 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	14 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1054_update_start_
      -- 
    outputPort_1_Daemon_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(9) & outputPort_1_Daemon_CP_2424_elements(176) & outputPort_1_Daemon_CP_2424_elements(179);
      gj_outputPort_1_Daemon_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	11 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1054_sample_start__ps
      -- 
    outputPort_1_Daemon_CP_2424_elements(58) <= outputPort_1_Daemon_CP_2424_elements(11);
    -- CP-element group 59:  join  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	12 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1054_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(59) is bound as output of CP function.
    -- CP-element group 60:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	14 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1054_update_start__ps
      -- 
    outputPort_1_Daemon_CP_2424_elements(60) <= outputPort_1_Daemon_CP_2424_elements(14);
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	178 
    -- CP-element group 61: 	174 
    -- CP-element group 61: 	15 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1054_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1054_update_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(61) is bound as output of CP function.
    -- CP-element group 62:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	7 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1054_loopback_trigger
      -- 
    outputPort_1_Daemon_CP_2424_elements(62) <= outputPort_1_Daemon_CP_2424_elements(7);
    -- CP-element group 63:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1054_loopback_sample_req
      -- CP-element group 63: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1054_loopback_sample_req_ps
      -- 
    phi_stmt_1054_loopback_sample_req_2552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1054_loopback_sample_req_2552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(63), ack => phi_stmt_1054_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(63) is bound as output of CP function.
    -- CP-element group 64:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	8 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1054_entry_trigger
      -- 
    outputPort_1_Daemon_CP_2424_elements(64) <= outputPort_1_Daemon_CP_2424_elements(8);
    -- CP-element group 65:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1054_entry_sample_req
      -- CP-element group 65: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1054_entry_sample_req_ps
      -- 
    phi_stmt_1054_entry_sample_req_2555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1054_entry_sample_req_2555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(65), ack => phi_stmt_1054_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(65) is bound as output of CP function.
    -- CP-element group 66:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1054_phi_mux_ack
      -- CP-element group 66: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1054_phi_mux_ack_ps
      -- 
    phi_stmt_1054_phi_mux_ack_2558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1054_ack_0, ack => outputPort_1_Daemon_CP_2424_elements(66)); -- 
    -- CP-element group 67:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1056_sample_start__ps
      -- CP-element group 67: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1056_sample_completed__ps
      -- CP-element group 67: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1056_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1056_sample_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1056_update_start__ps
      -- CP-element group 68: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1056_update_start_
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	70 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1056_update_completed__ps
      -- 
    outputPort_1_Daemon_CP_2424_elements(69) <= outputPort_1_Daemon_CP_2424_elements(70);
    -- CP-element group 70:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	69 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1056_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(70) is a control-delay.
    cp_element_70_delay: control_delay_element  generic map(name => " 70_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_2424_elements(68), ack => outputPort_1_Daemon_CP_2424_elements(70), clk => clk, reset =>reset);
    -- CP-element group 71:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_2_1_1058_sample_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(71) is bound as output of CP function.
    -- CP-element group 72:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_2_1_1058_update_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(72) is bound as output of CP function.
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: marked-predecessors 
    -- CP-element group 73: 	76 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_2_1_1058_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_2_1_1058_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_2_1_1058_Sample/rr
      -- 
    rr_2579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(73), ack => RPIPE_noblock_obuf_2_1_1058_inst_req_0); -- 
    outputPort_1_Daemon_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(71) & outputPort_1_Daemon_CP_2424_elements(76);
      gj_outputPort_1_Daemon_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: 	75 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_2_1_1058_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_2_1_1058_Update/cr
      -- CP-element group 74: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_2_1_1058_update_start_
      -- 
    cr_2584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(74), ack => RPIPE_noblock_obuf_2_1_1058_inst_req_1); -- 
    outputPort_1_Daemon_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(72) & outputPort_1_Daemon_CP_2424_elements(75);
      gj_outputPort_1_Daemon_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	74 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_2_1_1058_sample_completed__ps
      -- CP-element group 75: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_2_1_1058_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_2_1_1058_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_2_1_1058_Sample/ra
      -- 
    ra_2580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_1_1058_inst_ack_0, ack => outputPort_1_Daemon_CP_2424_elements(75)); -- 
    -- CP-element group 76:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: marked-successors 
    -- CP-element group 76: 	73 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_2_1_1058_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_2_1_1058_Update/ca
      -- CP-element group 76: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_2_1_1058_update_completed__ps
      -- CP-element group 76: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_2_1_1058_Update/$exit
      -- 
    ca_2585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_1_1058_inst_ack_1, ack => outputPort_1_Daemon_CP_2424_elements(76)); -- 
    -- CP-element group 77:  join  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	9 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	12 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	11 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1059_sample_start_
      -- 
    outputPort_1_Daemon_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(9) & outputPort_1_Daemon_CP_2424_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  join  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	9 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	176 
    -- CP-element group 78: 	179 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	14 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1059_update_start_
      -- 
    outputPort_1_Daemon_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(9) & outputPort_1_Daemon_CP_2424_elements(176) & outputPort_1_Daemon_CP_2424_elements(179);
      gj_outputPort_1_Daemon_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	11 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1059_sample_start__ps
      -- 
    outputPort_1_Daemon_CP_2424_elements(79) <= outputPort_1_Daemon_CP_2424_elements(11);
    -- CP-element group 80:  join  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	12 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1059_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(80) is bound as output of CP function.
    -- CP-element group 81:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	14 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1059_update_start__ps
      -- 
    outputPort_1_Daemon_CP_2424_elements(81) <= outputPort_1_Daemon_CP_2424_elements(14);
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	178 
    -- CP-element group 82: 	174 
    -- CP-element group 82: 	15 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1059_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1059_update_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(82) is bound as output of CP function.
    -- CP-element group 83:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	7 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1059_loopback_trigger
      -- 
    outputPort_1_Daemon_CP_2424_elements(83) <= outputPort_1_Daemon_CP_2424_elements(7);
    -- CP-element group 84:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1059_loopback_sample_req
      -- CP-element group 84: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1059_loopback_sample_req_ps
      -- 
    phi_stmt_1059_loopback_sample_req_2596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1059_loopback_sample_req_2596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(84), ack => phi_stmt_1059_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(84) is bound as output of CP function.
    -- CP-element group 85:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	8 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1059_entry_trigger
      -- 
    outputPort_1_Daemon_CP_2424_elements(85) <= outputPort_1_Daemon_CP_2424_elements(8);
    -- CP-element group 86:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1059_entry_sample_req
      -- CP-element group 86: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1059_entry_sample_req_ps
      -- 
    phi_stmt_1059_entry_sample_req_2599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1059_entry_sample_req_2599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(86), ack => phi_stmt_1059_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(86) is bound as output of CP function.
    -- CP-element group 87:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1059_phi_mux_ack_ps
      -- CP-element group 87: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1059_phi_mux_ack
      -- 
    phi_stmt_1059_phi_mux_ack_2602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1059_ack_0, ack => outputPort_1_Daemon_CP_2424_elements(87)); -- 
    -- CP-element group 88:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (4) 
      -- CP-element group 88: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1061_sample_start__ps
      -- CP-element group 88: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1061_sample_completed__ps
      -- CP-element group 88: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1061_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1061_sample_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1061_update_start__ps
      -- CP-element group 89: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1061_update_start_
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(89) is bound as output of CP function.
    -- CP-element group 90:  join  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	91 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1061_update_completed__ps
      -- 
    outputPort_1_Daemon_CP_2424_elements(90) <= outputPort_1_Daemon_CP_2424_elements(91);
    -- CP-element group 91:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	90 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1061_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(91) is a control-delay.
    cp_element_91_delay: control_delay_element  generic map(name => " 91_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_2424_elements(89), ack => outputPort_1_Daemon_CP_2424_elements(91), clk => clk, reset =>reset);
    -- CP-element group 92:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_3_1_1063_sample_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(92) is bound as output of CP function.
    -- CP-element group 93:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_3_1_1063_update_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(93) is bound as output of CP function.
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	97 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_3_1_1063_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_3_1_1063_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_3_1_1063_Sample/rr
      -- 
    rr_2623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(94), ack => RPIPE_noblock_obuf_3_1_1063_inst_req_0); -- 
    outputPort_1_Daemon_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(92) & outputPort_1_Daemon_CP_2424_elements(97);
      gj_outputPort_1_Daemon_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_3_1_1063_Update/$entry
      -- CP-element group 95: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_3_1_1063_Update/cr
      -- CP-element group 95: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_3_1_1063_update_start_
      -- 
    cr_2628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(95), ack => RPIPE_noblock_obuf_3_1_1063_inst_req_1); -- 
    outputPort_1_Daemon_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(96) & outputPort_1_Daemon_CP_2424_elements(93);
      gj_outputPort_1_Daemon_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	95 
    -- CP-element group 96:  members (4) 
      -- CP-element group 96: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_3_1_1063_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_3_1_1063_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_3_1_1063_Sample/ra
      -- CP-element group 96: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_3_1_1063_sample_completed__ps
      -- 
    ra_2624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_1_1063_inst_ack_0, ack => outputPort_1_Daemon_CP_2424_elements(96)); -- 
    -- CP-element group 97:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: marked-successors 
    -- CP-element group 97: 	94 
    -- CP-element group 97:  members (4) 
      -- CP-element group 97: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_3_1_1063_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_3_1_1063_Update/ca
      -- CP-element group 97: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_3_1_1063_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_3_1_1063_update_completed__ps
      -- 
    ca_2629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_1_1063_inst_ack_1, ack => outputPort_1_Daemon_CP_2424_elements(97)); -- 
    -- CP-element group 98:  join  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	9 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	12 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	11 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1064_sample_start_
      -- 
    outputPort_1_Daemon_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(9) & outputPort_1_Daemon_CP_2424_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  join  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	9 
    -- CP-element group 99: marked-predecessors 
    -- CP-element group 99: 	176 
    -- CP-element group 99: 	179 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	14 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1064_update_start_
      -- 
    outputPort_1_Daemon_cp_element_group_99: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_99"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(9) & outputPort_1_Daemon_CP_2424_elements(176) & outputPort_1_Daemon_CP_2424_elements(179);
      gj_outputPort_1_Daemon_cp_element_group_99 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(99), clk => clk, reset => reset); --
    end block;
    -- CP-element group 100:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	11 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1064_sample_start__ps
      -- 
    outputPort_1_Daemon_CP_2424_elements(100) <= outputPort_1_Daemon_CP_2424_elements(11);
    -- CP-element group 101:  join  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	12 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1064_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(101) is bound as output of CP function.
    -- CP-element group 102:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	14 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1064_update_start__ps
      -- 
    outputPort_1_Daemon_CP_2424_elements(102) <= outputPort_1_Daemon_CP_2424_elements(14);
    -- CP-element group 103:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	178 
    -- CP-element group 103: 	174 
    -- CP-element group 103: 	15 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1064_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1064_update_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(103) is bound as output of CP function.
    -- CP-element group 104:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	7 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1064_loopback_trigger
      -- 
    outputPort_1_Daemon_CP_2424_elements(104) <= outputPort_1_Daemon_CP_2424_elements(7);
    -- CP-element group 105:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1064_loopback_sample_req
      -- CP-element group 105: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1064_loopback_sample_req_ps
      -- 
    phi_stmt_1064_loopback_sample_req_2640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1064_loopback_sample_req_2640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(105), ack => phi_stmt_1064_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(105) is bound as output of CP function.
    -- CP-element group 106:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	8 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1064_entry_trigger
      -- 
    outputPort_1_Daemon_CP_2424_elements(106) <= outputPort_1_Daemon_CP_2424_elements(8);
    -- CP-element group 107:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1064_entry_sample_req
      -- CP-element group 107: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1064_entry_sample_req_ps
      -- 
    phi_stmt_1064_entry_sample_req_2643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1064_entry_sample_req_2643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(107), ack => phi_stmt_1064_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(107) is bound as output of CP function.
    -- CP-element group 108:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1064_phi_mux_ack
      -- CP-element group 108: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1064_phi_mux_ack_ps
      -- 
    phi_stmt_1064_phi_mux_ack_2646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1064_ack_0, ack => outputPort_1_Daemon_CP_2424_elements(108)); -- 
    -- CP-element group 109:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (4) 
      -- CP-element group 109: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1066_sample_start__ps
      -- CP-element group 109: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1066_sample_completed__ps
      -- CP-element group 109: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1066_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1066_sample_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(109) is bound as output of CP function.
    -- CP-element group 110:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1066_update_start__ps
      -- CP-element group 110: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1066_update_start_
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(110) is bound as output of CP function.
    -- CP-element group 111:  join  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1066_update_completed__ps
      -- 
    outputPort_1_Daemon_CP_2424_elements(111) <= outputPort_1_Daemon_CP_2424_elements(112);
    -- CP-element group 112:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	111 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_33_1066_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(112) is a control-delay.
    cp_element_112_delay: control_delay_element  generic map(name => " 112_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_2424_elements(110), ack => outputPort_1_Daemon_CP_2424_elements(112), clk => clk, reset =>reset);
    -- CP-element group 113:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_4_1_1068_sample_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(113) is bound as output of CP function.
    -- CP-element group 114:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_4_1_1068_update_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(114) is bound as output of CP function.
    -- CP-element group 115:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: marked-predecessors 
    -- CP-element group 115: 	118 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_4_1_1068_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_4_1_1068_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_4_1_1068_Sample/rr
      -- 
    rr_2667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(115), ack => RPIPE_noblock_obuf_4_1_1068_inst_req_0); -- 
    outputPort_1_Daemon_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(113) & outputPort_1_Daemon_CP_2424_elements(118);
      gj_outputPort_1_Daemon_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	117 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_4_1_1068_update_start_
      -- CP-element group 116: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_4_1_1068_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_4_1_1068_Update/cr
      -- 
    cr_2672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(116), ack => RPIPE_noblock_obuf_4_1_1068_inst_req_1); -- 
    outputPort_1_Daemon_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(117) & outputPort_1_Daemon_CP_2424_elements(114);
      gj_outputPort_1_Daemon_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	116 
    -- CP-element group 117:  members (4) 
      -- CP-element group 117: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_4_1_1068_sample_completed__ps
      -- CP-element group 117: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_4_1_1068_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_4_1_1068_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_4_1_1068_Sample/ra
      -- 
    ra_2668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_1_1068_inst_ack_0, ack => outputPort_1_Daemon_CP_2424_elements(117)); -- 
    -- CP-element group 118:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: marked-successors 
    -- CP-element group 118: 	115 
    -- CP-element group 118:  members (4) 
      -- CP-element group 118: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_4_1_1068_update_completed__ps
      -- CP-element group 118: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_4_1_1068_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_4_1_1068_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/RPIPE_noblock_obuf_4_1_1068_Update/ca
      -- 
    ca_2673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_1_1068_inst_ack_1, ack => outputPort_1_Daemon_CP_2424_elements(118)); -- 
    -- CP-element group 119:  join  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	9 
    -- CP-element group 119: marked-predecessors 
    -- CP-element group 119: 	12 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	11 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1069_sample_start_
      -- 
    outputPort_1_Daemon_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(9) & outputPort_1_Daemon_CP_2424_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  join  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	9 
    -- CP-element group 120: marked-predecessors 
    -- CP-element group 120: 	176 
    -- CP-element group 120: 	179 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	14 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1069_update_start_
      -- 
    outputPort_1_Daemon_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(9) & outputPort_1_Daemon_CP_2424_elements(176) & outputPort_1_Daemon_CP_2424_elements(179);
      gj_outputPort_1_Daemon_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  join  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	12 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1069_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(121) is bound as output of CP function.
    -- CP-element group 122:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	178 
    -- CP-element group 122: 	174 
    -- CP-element group 122: 	15 
    -- CP-element group 122:  members (2) 
      -- CP-element group 122: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1069_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1069_update_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(122) is bound as output of CP function.
    -- CP-element group 123:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	7 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1069_loopback_trigger
      -- 
    outputPort_1_Daemon_CP_2424_elements(123) <= outputPort_1_Daemon_CP_2424_elements(7);
    -- CP-element group 124:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (2) 
      -- CP-element group 124: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1069_loopback_sample_req
      -- CP-element group 124: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1069_loopback_sample_req_ps
      -- 
    phi_stmt_1069_loopback_sample_req_2684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1069_loopback_sample_req_2684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(124), ack => phi_stmt_1069_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(124) is bound as output of CP function.
    -- CP-element group 125:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	8 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1069_entry_trigger
      -- 
    outputPort_1_Daemon_CP_2424_elements(125) <= outputPort_1_Daemon_CP_2424_elements(8);
    -- CP-element group 126:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1069_entry_sample_req
      -- CP-element group 126: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1069_entry_sample_req_ps
      -- 
    phi_stmt_1069_entry_sample_req_2687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1069_entry_sample_req_2687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(126), ack => phi_stmt_1069_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(126) is bound as output of CP function.
    -- CP-element group 127:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1069_phi_mux_ack
      -- CP-element group 127: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1069_phi_mux_ack_ps
      -- 
    phi_stmt_1069_phi_mux_ack_2690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1069_ack_0, ack => outputPort_1_Daemon_CP_2424_elements(127)); -- 
    -- CP-element group 128:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (4) 
      -- CP-element group 128: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_3_1071_sample_start__ps
      -- CP-element group 128: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_3_1071_sample_completed__ps
      -- CP-element group 128: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_3_1071_sample_start_
      -- CP-element group 128: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_3_1071_sample_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(128) is bound as output of CP function.
    -- CP-element group 129:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	131 
    -- CP-element group 129:  members (2) 
      -- CP-element group 129: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_3_1071_update_start__ps
      -- CP-element group 129: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_3_1071_update_start_
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(129) is bound as output of CP function.
    -- CP-element group 130:  join  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: successors 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_3_1071_update_completed__ps
      -- 
    outputPort_1_Daemon_CP_2424_elements(130) <= outputPort_1_Daemon_CP_2424_elements(131);
    -- CP-element group 131:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	129 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	130 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_3_1071_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(131) is a control-delay.
    cp_element_131_delay: control_delay_element  generic map(name => " 131_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_2424_elements(129), ack => outputPort_1_Daemon_CP_2424_elements(131), clk => clk, reset =>reset);
    -- CP-element group 132:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (4) 
      -- CP-element group 132: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_1072_sample_start__ps
      -- CP-element group 132: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_1072_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_1072_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_1072_Sample/req
      -- 
    req_2711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(132), ack => next_active_packet_1179_1072_buf_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(132) is bound as output of CP function.
    -- CP-element group 133:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	135 
    -- CP-element group 133:  members (4) 
      -- CP-element group 133: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_1072_update_start__ps
      -- CP-element group 133: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_1072_update_start_
      -- CP-element group 133: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_1072_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_1072_Update/req
      -- 
    req_2716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(133), ack => next_active_packet_1179_1072_buf_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(133) is bound as output of CP function.
    -- CP-element group 134:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134:  members (4) 
      -- CP-element group 134: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_1072_sample_completed__ps
      -- CP-element group 134: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_1072_sample_completed_
      -- CP-element group 134: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_1072_Sample/$exit
      -- CP-element group 134: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_1072_Sample/ack
      -- 
    ack_2712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_1179_1072_buf_ack_0, ack => outputPort_1_Daemon_CP_2424_elements(134)); -- 
    -- CP-element group 135:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	133 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (4) 
      -- CP-element group 135: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_1072_update_completed__ps
      -- CP-element group 135: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_1072_update_completed_
      -- CP-element group 135: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_1072_Update/$exit
      -- CP-element group 135: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_1072_Update/ack
      -- 
    ack_2717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_1179_1072_buf_ack_1, ack => outputPort_1_Daemon_CP_2424_elements(135)); -- 
    -- CP-element group 136:  join  transition  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	9 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	12 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	11 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1073_sample_start_
      -- 
    outputPort_1_Daemon_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(9) & outputPort_1_Daemon_CP_2424_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  join  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	9 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	141 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	14 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1073_update_start_
      -- 
    outputPort_1_Daemon_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(9) & outputPort_1_Daemon_CP_2424_elements(141);
      gj_outputPort_1_Daemon_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	11 
    -- CP-element group 138: successors 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1073_sample_start__ps
      -- 
    outputPort_1_Daemon_CP_2424_elements(138) <= outputPort_1_Daemon_CP_2424_elements(11);
    -- CP-element group 139:  join  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	12 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1073_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(139) is bound as output of CP function.
    -- CP-element group 140:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	14 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (1) 
      -- CP-element group 140: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1073_update_start__ps
      -- 
    outputPort_1_Daemon_CP_2424_elements(140) <= outputPort_1_Daemon_CP_2424_elements(14);
    -- CP-element group 141:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	15 
    -- CP-element group 141: marked-successors 
    -- CP-element group 141: 	137 
    -- CP-element group 141:  members (2) 
      -- CP-element group 141: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1073_update_completed_
      -- CP-element group 141: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1073_update_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(141) is bound as output of CP function.
    -- CP-element group 142:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	7 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (1) 
      -- CP-element group 142: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1073_loopback_trigger
      -- 
    outputPort_1_Daemon_CP_2424_elements(142) <= outputPort_1_Daemon_CP_2424_elements(7);
    -- CP-element group 143:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (2) 
      -- CP-element group 143: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1073_loopback_sample_req
      -- CP-element group 143: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1073_loopback_sample_req_ps
      -- 
    phi_stmt_1073_loopback_sample_req_2728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1073_loopback_sample_req_2728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(143), ack => phi_stmt_1073_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(143) is bound as output of CP function.
    -- CP-element group 144:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	8 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (1) 
      -- CP-element group 144: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1073_entry_trigger
      -- 
    outputPort_1_Daemon_CP_2424_elements(144) <= outputPort_1_Daemon_CP_2424_elements(8);
    -- CP-element group 145:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1073_entry_sample_req
      -- CP-element group 145: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1073_entry_sample_req_ps
      -- 
    phi_stmt_1073_entry_sample_req_2731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1073_entry_sample_req_2731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(145), ack => phi_stmt_1073_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(145) is bound as output of CP function.
    -- CP-element group 146:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (2) 
      -- CP-element group 146: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1073_phi_mux_ack
      -- CP-element group 146: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1073_phi_mux_ack_ps
      -- 
    phi_stmt_1073_phi_mux_ack_2734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1073_ack_0, ack => outputPort_1_Daemon_CP_2424_elements(146)); -- 
    -- CP-element group 147:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (4) 
      -- CP-element group 147: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_8_1075_sample_start__ps
      -- CP-element group 147: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_8_1075_sample_completed__ps
      -- CP-element group 147: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_8_1075_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_8_1075_sample_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(147) is bound as output of CP function.
    -- CP-element group 148:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	150 
    -- CP-element group 148:  members (2) 
      -- CP-element group 148: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_8_1075_update_start__ps
      -- CP-element group 148: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_8_1075_update_start_
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(148) is bound as output of CP function.
    -- CP-element group 149:  join  transition  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	150 
    -- CP-element group 149: successors 
    -- CP-element group 149:  members (1) 
      -- CP-element group 149: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_8_1075_update_completed__ps
      -- 
    outputPort_1_Daemon_CP_2424_elements(149) <= outputPort_1_Daemon_CP_2424_elements(150);
    -- CP-element group 150:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	148 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	149 
    -- CP-element group 150:  members (1) 
      -- CP-element group 150: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_8_1075_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(150) is a control-delay.
    cp_element_150_delay: control_delay_element  generic map(name => " 150_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_2424_elements(148), ack => outputPort_1_Daemon_CP_2424_elements(150), clk => clk, reset =>reset);
    -- CP-element group 151:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (4) 
      -- CP-element group 151: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_length_1076_sample_start__ps
      -- CP-element group 151: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_length_1076_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_length_1076_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_length_1076_Sample/req
      -- 
    req_2755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(151), ack => next_active_packet_length_1224_1076_buf_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(151) is bound as output of CP function.
    -- CP-element group 152:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (4) 
      -- CP-element group 152: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_length_1076_update_start__ps
      -- CP-element group 152: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_length_1076_update_start_
      -- CP-element group 152: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_length_1076_Update/$entry
      -- CP-element group 152: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_length_1076_Update/req
      -- 
    req_2760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(152), ack => next_active_packet_length_1224_1076_buf_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(152) is bound as output of CP function.
    -- CP-element group 153:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (4) 
      -- CP-element group 153: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_length_1076_sample_completed__ps
      -- CP-element group 153: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_length_1076_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_length_1076_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_length_1076_Sample/ack
      -- 
    ack_2756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_length_1224_1076_buf_ack_0, ack => outputPort_1_Daemon_CP_2424_elements(153)); -- 
    -- CP-element group 154:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	152 
    -- CP-element group 154: successors 
    -- CP-element group 154:  members (4) 
      -- CP-element group 154: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_length_1076_update_completed__ps
      -- CP-element group 154: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_length_1076_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_length_1076_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_active_packet_length_1076_Update/ack
      -- 
    ack_2761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_length_1224_1076_buf_ack_1, ack => outputPort_1_Daemon_CP_2424_elements(154)); -- 
    -- CP-element group 155:  join  transition  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	9 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	12 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	11 
    -- CP-element group 155:  members (1) 
      -- CP-element group 155: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1077_sample_start_
      -- 
    outputPort_1_Daemon_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(9) & outputPort_1_Daemon_CP_2424_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  join  transition  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	9 
    -- CP-element group 156: marked-predecessors 
    -- CP-element group 156: 	176 
    -- CP-element group 156: 	179 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	14 
    -- CP-element group 156:  members (1) 
      -- CP-element group 156: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1077_update_start_
      -- 
    outputPort_1_Daemon_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(9) & outputPort_1_Daemon_CP_2424_elements(176) & outputPort_1_Daemon_CP_2424_elements(179);
      gj_outputPort_1_Daemon_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	11 
    -- CP-element group 157: successors 
    -- CP-element group 157:  members (1) 
      -- CP-element group 157: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1077_sample_start__ps
      -- 
    outputPort_1_Daemon_CP_2424_elements(157) <= outputPort_1_Daemon_CP_2424_elements(11);
    -- CP-element group 158:  join  transition  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	12 
    -- CP-element group 158:  members (1) 
      -- CP-element group 158: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1077_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(158) is bound as output of CP function.
    -- CP-element group 159:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	14 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (1) 
      -- CP-element group 159: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1077_update_start__ps
      -- 
    outputPort_1_Daemon_CP_2424_elements(159) <= outputPort_1_Daemon_CP_2424_elements(14);
    -- CP-element group 160:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	178 
    -- CP-element group 160: 	174 
    -- CP-element group 160: 	15 
    -- CP-element group 160:  members (2) 
      -- CP-element group 160: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1077_update_completed_
      -- CP-element group 160: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1077_update_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(160) is bound as output of CP function.
    -- CP-element group 161:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	7 
    -- CP-element group 161: successors 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1077_loopback_trigger
      -- 
    outputPort_1_Daemon_CP_2424_elements(161) <= outputPort_1_Daemon_CP_2424_elements(7);
    -- CP-element group 162:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (2) 
      -- CP-element group 162: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1077_loopback_sample_req
      -- CP-element group 162: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1077_loopback_sample_req_ps
      -- 
    phi_stmt_1077_loopback_sample_req_2772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1077_loopback_sample_req_2772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(162), ack => phi_stmt_1077_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(162) is bound as output of CP function.
    -- CP-element group 163:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	8 
    -- CP-element group 163: successors 
    -- CP-element group 163:  members (1) 
      -- CP-element group 163: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1077_entry_trigger
      -- 
    outputPort_1_Daemon_CP_2424_elements(163) <= outputPort_1_Daemon_CP_2424_elements(8);
    -- CP-element group 164:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (2) 
      -- CP-element group 164: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1077_entry_sample_req
      -- CP-element group 164: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1077_entry_sample_req_ps
      -- 
    phi_stmt_1077_entry_sample_req_2775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1077_entry_sample_req_2775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(164), ack => phi_stmt_1077_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(164) is bound as output of CP function.
    -- CP-element group 165:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: successors 
    -- CP-element group 165:  members (2) 
      -- CP-element group 165: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1077_phi_mux_ack
      -- CP-element group 165: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/phi_stmt_1077_phi_mux_ack_ps
      -- 
    phi_stmt_1077_phi_mux_ack_2778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1077_ack_0, ack => outputPort_1_Daemon_CP_2424_elements(165)); -- 
    -- CP-element group 166:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: successors 
    -- CP-element group 166:  members (4) 
      -- CP-element group 166: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_2_1079_sample_start__ps
      -- CP-element group 166: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_2_1079_sample_completed__ps
      -- CP-element group 166: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_2_1079_sample_start_
      -- CP-element group 166: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_2_1079_sample_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(166) is bound as output of CP function.
    -- CP-element group 167:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (2) 
      -- CP-element group 167: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_2_1079_update_start__ps
      -- CP-element group 167: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_2_1079_update_start_
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(167) is bound as output of CP function.
    -- CP-element group 168:  join  transition  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	169 
    -- CP-element group 168: successors 
    -- CP-element group 168:  members (1) 
      -- CP-element group 168: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_2_1079_update_completed__ps
      -- 
    outputPort_1_Daemon_CP_2424_elements(168) <= outputPort_1_Daemon_CP_2424_elements(169);
    -- CP-element group 169:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	168 
    -- CP-element group 169:  members (1) 
      -- CP-element group 169: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_ZERO_2_1079_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(169) is a control-delay.
    cp_element_169_delay: control_delay_element  generic map(name => " 169_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_2424_elements(167), ack => outputPort_1_Daemon_CP_2424_elements(169), clk => clk, reset =>reset);
    -- CP-element group 170:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	172 
    -- CP-element group 170:  members (4) 
      -- CP-element group 170: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_priority_index_1080_sample_start__ps
      -- CP-element group 170: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_priority_index_1080_sample_start_
      -- CP-element group 170: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_priority_index_1080_Sample/$entry
      -- CP-element group 170: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_priority_index_1080_Sample/req
      -- 
    req_2799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(170), ack => next_priority_index_1179_1080_buf_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(170) is bound as output of CP function.
    -- CP-element group 171:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (4) 
      -- CP-element group 171: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_priority_index_1080_update_start__ps
      -- CP-element group 171: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_priority_index_1080_update_start_
      -- CP-element group 171: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_priority_index_1080_Update/$entry
      -- CP-element group 171: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_priority_index_1080_Update/req
      -- 
    req_2804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(171), ack => next_priority_index_1179_1080_buf_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(171) is bound as output of CP function.
    -- CP-element group 172:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	170 
    -- CP-element group 172: successors 
    -- CP-element group 172:  members (4) 
      -- CP-element group 172: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_priority_index_1080_sample_completed__ps
      -- CP-element group 172: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_priority_index_1080_sample_completed_
      -- CP-element group 172: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_priority_index_1080_Sample/$exit
      -- CP-element group 172: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_priority_index_1080_Sample/ack
      -- 
    ack_2800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_priority_index_1179_1080_buf_ack_0, ack => outputPort_1_Daemon_CP_2424_elements(172)); -- 
    -- CP-element group 173:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: successors 
    -- CP-element group 173:  members (4) 
      -- CP-element group 173: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_priority_index_1080_update_completed__ps
      -- CP-element group 173: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_priority_index_1080_update_completed_
      -- CP-element group 173: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_priority_index_1080_Update/$exit
      -- CP-element group 173: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/R_next_priority_index_1080_Update/ack
      -- 
    ack_2805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_priority_index_1179_1080_buf_ack_1, ack => outputPort_1_Daemon_CP_2424_elements(173)); -- 
    -- CP-element group 174:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	122 
    -- CP-element group 174: 	160 
    -- CP-element group 174: 	21 
    -- CP-element group 174: 	40 
    -- CP-element group 174: 	103 
    -- CP-element group 174: 	61 
    -- CP-element group 174: 	82 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	176 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/call_stmt_1108_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/call_stmt_1108_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/call_stmt_1108_Sample/crr
      -- 
    crr_2814_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2814_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(174), ack => call_stmt_1108_call_req_0); -- 
    outputPort_1_Daemon_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(122) & outputPort_1_Daemon_CP_2424_elements(160) & outputPort_1_Daemon_CP_2424_elements(21) & outputPort_1_Daemon_CP_2424_elements(40) & outputPort_1_Daemon_CP_2424_elements(103) & outputPort_1_Daemon_CP_2424_elements(61) & outputPort_1_Daemon_CP_2424_elements(82);
      gj_outputPort_1_Daemon_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: marked-predecessors 
    -- CP-element group 175: 	177 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	177 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/call_stmt_1108_update_start_
      -- CP-element group 175: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/call_stmt_1108_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/call_stmt_1108_Update/ccr
      -- 
    ccr_2819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(175), ack => call_stmt_1108_call_req_1); -- 
    outputPort_1_Daemon_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= outputPort_1_Daemon_CP_2424_elements(177);
      gj_outputPort_1_Daemon_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	174 
    -- CP-element group 176: successors 
    -- CP-element group 176: marked-successors 
    -- CP-element group 176: 	99 
    -- CP-element group 176: 	120 
    -- CP-element group 176: 	156 
    -- CP-element group 176: 	17 
    -- CP-element group 176: 	36 
    -- CP-element group 176: 	57 
    -- CP-element group 176: 	78 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/call_stmt_1108_sample_completed_
      -- CP-element group 176: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/call_stmt_1108_Sample/$exit
      -- CP-element group 176: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/call_stmt_1108_Sample/cra
      -- 
    cra_2815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1108_call_ack_0, ack => outputPort_1_Daemon_CP_2424_elements(176)); -- 
    -- CP-element group 177:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	182 
    -- CP-element group 177: marked-successors 
    -- CP-element group 177: 	175 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/call_stmt_1108_update_completed_
      -- CP-element group 177: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/call_stmt_1108_Update/$exit
      -- CP-element group 177: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/call_stmt_1108_Update/cca
      -- 
    cca_2820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1108_call_ack_1, ack => outputPort_1_Daemon_CP_2424_elements(177)); -- 
    -- CP-element group 178:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	122 
    -- CP-element group 178: 	160 
    -- CP-element group 178: 	21 
    -- CP-element group 178: 	40 
    -- CP-element group 178: 	103 
    -- CP-element group 178: 	61 
    -- CP-element group 178: 	82 
    -- CP-element group 178: marked-predecessors 
    -- CP-element group 178: 	180 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/WPIPE_out_data_1_1333_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/WPIPE_out_data_1_1333_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/WPIPE_out_data_1_1333_Sample/req
      -- 
    req_2828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(178), ack => WPIPE_out_data_1_1333_inst_req_0); -- 
    outputPort_1_Daemon_cp_element_group_178: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_178"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(122) & outputPort_1_Daemon_CP_2424_elements(160) & outputPort_1_Daemon_CP_2424_elements(21) & outputPort_1_Daemon_CP_2424_elements(40) & outputPort_1_Daemon_CP_2424_elements(103) & outputPort_1_Daemon_CP_2424_elements(61) & outputPort_1_Daemon_CP_2424_elements(82) & outputPort_1_Daemon_CP_2424_elements(180);
      gj_outputPort_1_Daemon_cp_element_group_178 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(178), clk => clk, reset => reset); --
    end block;
    -- CP-element group 179:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179: marked-successors 
    -- CP-element group 179: 	99 
    -- CP-element group 179: 	120 
    -- CP-element group 179: 	156 
    -- CP-element group 179: 	17 
    -- CP-element group 179: 	36 
    -- CP-element group 179: 	57 
    -- CP-element group 179: 	78 
    -- CP-element group 179:  members (6) 
      -- CP-element group 179: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/WPIPE_out_data_1_1333_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/WPIPE_out_data_1_1333_update_start_
      -- CP-element group 179: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/WPIPE_out_data_1_1333_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/WPIPE_out_data_1_1333_Sample/ack
      -- CP-element group 179: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/WPIPE_out_data_1_1333_Update/$entry
      -- CP-element group 179: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/WPIPE_out_data_1_1333_Update/req
      -- 
    ack_2829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_1_1333_inst_ack_0, ack => outputPort_1_Daemon_CP_2424_elements(179)); -- 
    req_2833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_2424_elements(179), ack => WPIPE_out_data_1_1333_inst_req_1); -- 
    -- CP-element group 180:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	182 
    -- CP-element group 180: marked-successors 
    -- CP-element group 180: 	178 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/WPIPE_out_data_1_1333_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/WPIPE_out_data_1_1333_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/WPIPE_out_data_1_1333_Update/ack
      -- 
    ack_2834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_1_1333_inst_ack_1, ack => outputPort_1_Daemon_CP_2424_elements(180)); -- 
    -- CP-element group 181:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	9 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	10 
    -- CP-element group 181:  members (1) 
      -- CP-element group 181: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group outputPort_1_Daemon_CP_2424_elements(181) is a control-delay.
    cp_element_181_delay: control_delay_element  generic map(name => " 181_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_2424_elements(9), ack => outputPort_1_Daemon_CP_2424_elements(181), clk => clk, reset =>reset);
    -- CP-element group 182:  join  transition  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	177 
    -- CP-element group 182: 	180 
    -- CP-element group 182: 	12 
    -- CP-element group 182: 	13 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	6 
    -- CP-element group 182:  members (1) 
      -- CP-element group 182: 	 branch_block_stmt_1042/do_while_stmt_1043/do_while_stmt_1043_loop_body/$exit
      -- 
    outputPort_1_Daemon_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 7,2 => 7,3 => 7);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_2424_elements(177) & outputPort_1_Daemon_CP_2424_elements(180) & outputPort_1_Daemon_CP_2424_elements(12) & outputPort_1_Daemon_CP_2424_elements(13);
      gj_outputPort_1_Daemon_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  transition  input  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	5 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (2) 
      -- CP-element group 183: 	 branch_block_stmt_1042/do_while_stmt_1043/loop_exit/$exit
      -- CP-element group 183: 	 branch_block_stmt_1042/do_while_stmt_1043/loop_exit/ack
      -- 
    ack_2839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1043_branch_ack_0, ack => outputPort_1_Daemon_CP_2424_elements(183)); -- 
    -- CP-element group 184:  transition  input  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	5 
    -- CP-element group 184: successors 
    -- CP-element group 184:  members (2) 
      -- CP-element group 184: 	 branch_block_stmt_1042/do_while_stmt_1043/loop_taken/$exit
      -- CP-element group 184: 	 branch_block_stmt_1042/do_while_stmt_1043/loop_taken/ack
      -- 
    ack_2843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1043_branch_ack_1, ack => outputPort_1_Daemon_CP_2424_elements(184)); -- 
    -- CP-element group 185:  transition  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	3 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	1 
    -- CP-element group 185:  members (1) 
      -- CP-element group 185: 	 branch_block_stmt_1042/do_while_stmt_1043/$exit
      -- 
    outputPort_1_Daemon_CP_2424_elements(185) <= outputPort_1_Daemon_CP_2424_elements(3);
    outputPort_1_Daemon_do_while_stmt_1043_terminator_2844: loop_terminator -- 
      generic map (name => " outputPort_1_Daemon_do_while_stmt_1043_terminator_2844", max_iterations_in_flight =>7) 
      port map(loop_body_exit => outputPort_1_Daemon_CP_2424_elements(6),loop_continue => outputPort_1_Daemon_CP_2424_elements(184),loop_terminate => outputPort_1_Daemon_CP_2424_elements(183),loop_back => outputPort_1_Daemon_CP_2424_elements(4),loop_exit => outputPort_1_Daemon_CP_2424_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1045_phi_seq_2498_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_1_Daemon_CP_2424_elements(24);
      outputPort_1_Daemon_CP_2424_elements(27)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_1_Daemon_CP_2424_elements(27);
      outputPort_1_Daemon_CP_2424_elements(28)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_1_Daemon_CP_2424_elements(29);
      outputPort_1_Daemon_CP_2424_elements(25) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_1_Daemon_CP_2424_elements(22);
      outputPort_1_Daemon_CP_2424_elements(31)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_1_Daemon_CP_2424_elements(33);
      outputPort_1_Daemon_CP_2424_elements(32)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_1_Daemon_CP_2424_elements(34);
      outputPort_1_Daemon_CP_2424_elements(23) <= phi_mux_reqs(1);
      phi_stmt_1045_phi_seq_2498 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1045_phi_seq_2498") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_1_Daemon_CP_2424_elements(18), 
          phi_sample_ack => outputPort_1_Daemon_CP_2424_elements(19), 
          phi_update_req => outputPort_1_Daemon_CP_2424_elements(20), 
          phi_update_ack => outputPort_1_Daemon_CP_2424_elements(21), 
          phi_mux_ack => outputPort_1_Daemon_CP_2424_elements(26), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1049_phi_seq_2542_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_1_Daemon_CP_2424_elements(43);
      outputPort_1_Daemon_CP_2424_elements(46)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_1_Daemon_CP_2424_elements(46);
      outputPort_1_Daemon_CP_2424_elements(47)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_1_Daemon_CP_2424_elements(48);
      outputPort_1_Daemon_CP_2424_elements(44) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_1_Daemon_CP_2424_elements(41);
      outputPort_1_Daemon_CP_2424_elements(50)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_1_Daemon_CP_2424_elements(54);
      outputPort_1_Daemon_CP_2424_elements(51)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_1_Daemon_CP_2424_elements(55);
      outputPort_1_Daemon_CP_2424_elements(42) <= phi_mux_reqs(1);
      phi_stmt_1049_phi_seq_2542 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1049_phi_seq_2542") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_1_Daemon_CP_2424_elements(37), 
          phi_sample_ack => outputPort_1_Daemon_CP_2424_elements(38), 
          phi_update_req => outputPort_1_Daemon_CP_2424_elements(39), 
          phi_update_ack => outputPort_1_Daemon_CP_2424_elements(40), 
          phi_mux_ack => outputPort_1_Daemon_CP_2424_elements(45), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1054_phi_seq_2586_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_1_Daemon_CP_2424_elements(64);
      outputPort_1_Daemon_CP_2424_elements(67)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_1_Daemon_CP_2424_elements(67);
      outputPort_1_Daemon_CP_2424_elements(68)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_1_Daemon_CP_2424_elements(69);
      outputPort_1_Daemon_CP_2424_elements(65) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_1_Daemon_CP_2424_elements(62);
      outputPort_1_Daemon_CP_2424_elements(71)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_1_Daemon_CP_2424_elements(75);
      outputPort_1_Daemon_CP_2424_elements(72)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_1_Daemon_CP_2424_elements(76);
      outputPort_1_Daemon_CP_2424_elements(63) <= phi_mux_reqs(1);
      phi_stmt_1054_phi_seq_2586 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1054_phi_seq_2586") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_1_Daemon_CP_2424_elements(58), 
          phi_sample_ack => outputPort_1_Daemon_CP_2424_elements(59), 
          phi_update_req => outputPort_1_Daemon_CP_2424_elements(60), 
          phi_update_ack => outputPort_1_Daemon_CP_2424_elements(61), 
          phi_mux_ack => outputPort_1_Daemon_CP_2424_elements(66), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1059_phi_seq_2630_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_1_Daemon_CP_2424_elements(85);
      outputPort_1_Daemon_CP_2424_elements(88)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_1_Daemon_CP_2424_elements(88);
      outputPort_1_Daemon_CP_2424_elements(89)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_1_Daemon_CP_2424_elements(90);
      outputPort_1_Daemon_CP_2424_elements(86) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_1_Daemon_CP_2424_elements(83);
      outputPort_1_Daemon_CP_2424_elements(92)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_1_Daemon_CP_2424_elements(96);
      outputPort_1_Daemon_CP_2424_elements(93)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_1_Daemon_CP_2424_elements(97);
      outputPort_1_Daemon_CP_2424_elements(84) <= phi_mux_reqs(1);
      phi_stmt_1059_phi_seq_2630 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1059_phi_seq_2630") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_1_Daemon_CP_2424_elements(79), 
          phi_sample_ack => outputPort_1_Daemon_CP_2424_elements(80), 
          phi_update_req => outputPort_1_Daemon_CP_2424_elements(81), 
          phi_update_ack => outputPort_1_Daemon_CP_2424_elements(82), 
          phi_mux_ack => outputPort_1_Daemon_CP_2424_elements(87), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1064_phi_seq_2674_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_1_Daemon_CP_2424_elements(106);
      outputPort_1_Daemon_CP_2424_elements(109)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_1_Daemon_CP_2424_elements(109);
      outputPort_1_Daemon_CP_2424_elements(110)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_1_Daemon_CP_2424_elements(111);
      outputPort_1_Daemon_CP_2424_elements(107) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_1_Daemon_CP_2424_elements(104);
      outputPort_1_Daemon_CP_2424_elements(113)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_1_Daemon_CP_2424_elements(117);
      outputPort_1_Daemon_CP_2424_elements(114)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_1_Daemon_CP_2424_elements(118);
      outputPort_1_Daemon_CP_2424_elements(105) <= phi_mux_reqs(1);
      phi_stmt_1064_phi_seq_2674 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1064_phi_seq_2674") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_1_Daemon_CP_2424_elements(100), 
          phi_sample_ack => outputPort_1_Daemon_CP_2424_elements(101), 
          phi_update_req => outputPort_1_Daemon_CP_2424_elements(102), 
          phi_update_ack => outputPort_1_Daemon_CP_2424_elements(103), 
          phi_mux_ack => outputPort_1_Daemon_CP_2424_elements(108), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1069_phi_seq_2718_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_1_Daemon_CP_2424_elements(125);
      outputPort_1_Daemon_CP_2424_elements(128)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_1_Daemon_CP_2424_elements(128);
      outputPort_1_Daemon_CP_2424_elements(129)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_1_Daemon_CP_2424_elements(130);
      outputPort_1_Daemon_CP_2424_elements(126) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_1_Daemon_CP_2424_elements(123);
      outputPort_1_Daemon_CP_2424_elements(132)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_1_Daemon_CP_2424_elements(134);
      outputPort_1_Daemon_CP_2424_elements(133)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_1_Daemon_CP_2424_elements(135);
      outputPort_1_Daemon_CP_2424_elements(124) <= phi_mux_reqs(1);
      phi_stmt_1069_phi_seq_2718 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1069_phi_seq_2718") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_1_Daemon_CP_2424_elements(11), 
          phi_sample_ack => outputPort_1_Daemon_CP_2424_elements(121), 
          phi_update_req => outputPort_1_Daemon_CP_2424_elements(14), 
          phi_update_ack => outputPort_1_Daemon_CP_2424_elements(122), 
          phi_mux_ack => outputPort_1_Daemon_CP_2424_elements(127), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1073_phi_seq_2762_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_1_Daemon_CP_2424_elements(144);
      outputPort_1_Daemon_CP_2424_elements(147)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_1_Daemon_CP_2424_elements(147);
      outputPort_1_Daemon_CP_2424_elements(148)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_1_Daemon_CP_2424_elements(149);
      outputPort_1_Daemon_CP_2424_elements(145) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_1_Daemon_CP_2424_elements(142);
      outputPort_1_Daemon_CP_2424_elements(151)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_1_Daemon_CP_2424_elements(153);
      outputPort_1_Daemon_CP_2424_elements(152)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_1_Daemon_CP_2424_elements(154);
      outputPort_1_Daemon_CP_2424_elements(143) <= phi_mux_reqs(1);
      phi_stmt_1073_phi_seq_2762 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1073_phi_seq_2762") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_1_Daemon_CP_2424_elements(138), 
          phi_sample_ack => outputPort_1_Daemon_CP_2424_elements(139), 
          phi_update_req => outputPort_1_Daemon_CP_2424_elements(140), 
          phi_update_ack => outputPort_1_Daemon_CP_2424_elements(141), 
          phi_mux_ack => outputPort_1_Daemon_CP_2424_elements(146), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1077_phi_seq_2806_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_1_Daemon_CP_2424_elements(163);
      outputPort_1_Daemon_CP_2424_elements(166)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_1_Daemon_CP_2424_elements(166);
      outputPort_1_Daemon_CP_2424_elements(167)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_1_Daemon_CP_2424_elements(168);
      outputPort_1_Daemon_CP_2424_elements(164) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_1_Daemon_CP_2424_elements(161);
      outputPort_1_Daemon_CP_2424_elements(170)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_1_Daemon_CP_2424_elements(172);
      outputPort_1_Daemon_CP_2424_elements(171)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_1_Daemon_CP_2424_elements(173);
      outputPort_1_Daemon_CP_2424_elements(162) <= phi_mux_reqs(1);
      phi_stmt_1077_phi_seq_2806 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1077_phi_seq_2806") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_1_Daemon_CP_2424_elements(157), 
          phi_sample_ack => outputPort_1_Daemon_CP_2424_elements(158), 
          phi_update_req => outputPort_1_Daemon_CP_2424_elements(159), 
          phi_update_ack => outputPort_1_Daemon_CP_2424_elements(160), 
          phi_mux_ack => outputPort_1_Daemon_CP_2424_elements(165), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_2449_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= outputPort_1_Daemon_CP_2424_elements(7);
        preds(1)  <= outputPort_1_Daemon_CP_2424_elements(8);
        entry_tmerge_2449 : transition_merge -- 
          generic map(name => " entry_tmerge_2449")
          port map (preds => preds, symbol_out => outputPort_1_Daemon_CP_2424_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal EQ_u3_u1_1144_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1150_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1157_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1163_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1193_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1200_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1208_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1215_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1243_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1251_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1259_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1267_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1273_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1280_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1288_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1295_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1306_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1312_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1319_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1325_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_1186_wire : std_logic_vector(0 downto 0);
    signal MUX_1086_wire : std_logic_vector(7 downto 0);
    signal MUX_1090_wire : std_logic_vector(7 downto 0);
    signal MUX_1095_wire : std_logic_vector(7 downto 0);
    signal MUX_1099_wire : std_logic_vector(7 downto 0);
    signal MUX_1147_wire : std_logic_vector(0 downto 0);
    signal MUX_1153_wire : std_logic_vector(0 downto 0);
    signal MUX_1160_wire : std_logic_vector(0 downto 0);
    signal MUX_1166_wire : std_logic_vector(0 downto 0);
    signal MUX_1197_wire : std_logic_vector(7 downto 0);
    signal MUX_1204_wire : std_logic_vector(7 downto 0);
    signal MUX_1212_wire : std_logic_vector(7 downto 0);
    signal MUX_1219_wire : std_logic_vector(7 downto 0);
    signal MUX_1235_wire : std_logic_vector(7 downto 0);
    signal MUX_1277_wire : std_logic_vector(31 downto 0);
    signal MUX_1284_wire : std_logic_vector(31 downto 0);
    signal MUX_1292_wire : std_logic_vector(31 downto 0);
    signal MUX_1299_wire : std_logic_vector(31 downto 0);
    signal MUX_1309_wire : std_logic_vector(0 downto 0);
    signal MUX_1315_wire : std_logic_vector(0 downto 0);
    signal MUX_1322_wire : std_logic_vector(0 downto 0);
    signal MUX_1328_wire : std_logic_vector(0 downto 0);
    signal NEQ_u3_u1_1183_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1240_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1248_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1256_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1264_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1154_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1167_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1316_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1329_wire : std_logic_vector(0 downto 0);
    signal OR_u32_u32_1285_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_1300_wire : std_logic_vector(31 downto 0);
    signal OR_u8_u8_1091_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_1100_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_1205_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_1220_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_1221_wire : std_logic_vector(7 downto 0);
    signal RPIPE_noblock_obuf_1_1_1053_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_2_1_1058_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_3_1_1063_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_4_1_1068_wire : std_logic_vector(32 downto 0);
    signal R_ZERO_2_1079_wire_constant : std_logic_vector(1 downto 0);
    signal R_ZERO_33_1051_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1056_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1061_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1066_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_3_1071_wire_constant : std_logic_vector(2 downto 0);
    signal R_ZERO_8_1047_wire_constant : std_logic_vector(7 downto 0);
    signal R_ZERO_8_1075_wire_constant : std_logic_vector(7 downto 0);
    signal SUB_u8_u8_1229_wire : std_logic_vector(7 downto 0);
    signal SUB_u8_u8_1233_wire : std_logic_vector(7 downto 0);
    signal active_packet_1069 : std_logic_vector(2 downto 0);
    signal active_packet_length_1073 : std_logic_vector(7 downto 0);
    signal continue_1108 : std_logic_vector(0 downto 0);
    signal data_to_out_1302 : std_logic_vector(31 downto 0);
    signal down_counter_1045 : std_logic_vector(7 downto 0);
    signal konst_1084_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1085_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1088_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1089_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1093_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1094_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1097_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1098_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1104_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1111_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1116_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1121_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1126_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1143_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1146_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1149_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1152_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1156_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1159_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1162_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1165_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1182_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1185_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1192_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1196_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1199_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1203_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1207_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1211_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1214_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1218_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1228_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1232_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1242_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1250_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1258_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1266_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1272_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1276_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1279_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1283_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1287_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1291_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1294_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1298_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1305_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1308_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1311_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1314_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1318_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1321_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1324_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1327_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1346_wire_constant : std_logic_vector(0 downto 0);
    signal next_active_packet_1179 : std_logic_vector(2 downto 0);
    signal next_active_packet_1179_1072_buffered : std_logic_vector(2 downto 0);
    signal next_active_packet_length_1224 : std_logic_vector(7 downto 0);
    signal next_active_packet_length_1224_1076_buffered : std_logic_vector(7 downto 0);
    signal next_down_counter_1237 : std_logic_vector(7 downto 0);
    signal next_down_counter_1237_1048_buffered : std_logic_vector(7 downto 0);
    signal next_priority_index_1179 : std_logic_vector(1 downto 0);
    signal next_priority_index_1179_1080_buffered : std_logic_vector(1 downto 0);
    signal p1_valid_1113 : std_logic_vector(0 downto 0);
    signal p2_valid_1118 : std_logic_vector(0 downto 0);
    signal p3_valid_1123 : std_logic_vector(0 downto 0);
    signal p4_valid_1128 : std_logic_vector(0 downto 0);
    signal pkt_1_e_word_1049 : std_logic_vector(32 downto 0);
    signal pkt_2_e_word_1054 : std_logic_vector(32 downto 0);
    signal pkt_3_e_word_1059 : std_logic_vector(32 downto 0);
    signal pkt_4_e_word_1064 : std_logic_vector(32 downto 0);
    signal priority_index_1077 : std_logic_vector(1 downto 0);
    signal read_from_1_1245 : std_logic_vector(0 downto 0);
    signal read_from_2_1253 : std_logic_vector(0 downto 0);
    signal read_from_3_1261 : std_logic_vector(0 downto 0);
    signal read_from_4_1269 : std_logic_vector(0 downto 0);
    signal send_flag_1331 : std_logic_vector(0 downto 0);
    signal senderPort_1102 : std_logic_vector(7 downto 0);
    signal slice_1195_wire : std_logic_vector(7 downto 0);
    signal slice_1202_wire : std_logic_vector(7 downto 0);
    signal slice_1210_wire : std_logic_vector(7 downto 0);
    signal slice_1217_wire : std_logic_vector(7 downto 0);
    signal slice_1275_wire : std_logic_vector(31 downto 0);
    signal slice_1282_wire : std_logic_vector(31 downto 0);
    signal slice_1290_wire : std_logic_vector(31 downto 0);
    signal slice_1297_wire : std_logic_vector(31 downto 0);
    signal started_new_packet_1188 : std_logic_vector(0 downto 0);
    signal type_cast_1106_wire_constant : std_logic_vector(0 downto 0);
    signal valid_active_pkt_word_read_1169 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_ZERO_2_1079_wire_constant <= "00";
    R_ZERO_33_1051_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1056_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1061_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1066_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_3_1071_wire_constant <= "000";
    R_ZERO_8_1047_wire_constant <= "00000000";
    R_ZERO_8_1075_wire_constant <= "00000000";
    konst_1084_wire_constant <= "00000000";
    konst_1085_wire_constant <= "00000000";
    konst_1088_wire_constant <= "00000001";
    konst_1089_wire_constant <= "00000000";
    konst_1093_wire_constant <= "00000010";
    konst_1094_wire_constant <= "00000000";
    konst_1097_wire_constant <= "00000011";
    konst_1098_wire_constant <= "00000000";
    konst_1104_wire_constant <= "00000000";
    konst_1111_wire_constant <= "000000000000000000000000000100000";
    konst_1116_wire_constant <= "000000000000000000000000000100000";
    konst_1121_wire_constant <= "000000000000000000000000000100000";
    konst_1126_wire_constant <= "000000000000000000000000000100000";
    konst_1143_wire_constant <= "001";
    konst_1146_wire_constant <= "0";
    konst_1149_wire_constant <= "010";
    konst_1152_wire_constant <= "0";
    konst_1156_wire_constant <= "011";
    konst_1159_wire_constant <= "0";
    konst_1162_wire_constant <= "100";
    konst_1165_wire_constant <= "0";
    konst_1182_wire_constant <= "000";
    konst_1185_wire_constant <= "00000000";
    konst_1192_wire_constant <= "001";
    konst_1196_wire_constant <= "00000000";
    konst_1199_wire_constant <= "010";
    konst_1203_wire_constant <= "00000000";
    konst_1207_wire_constant <= "011";
    konst_1211_wire_constant <= "00000000";
    konst_1214_wire_constant <= "100";
    konst_1218_wire_constant <= "00000000";
    konst_1228_wire_constant <= "00000001";
    konst_1232_wire_constant <= "00000001";
    konst_1242_wire_constant <= "001";
    konst_1250_wire_constant <= "010";
    konst_1258_wire_constant <= "011";
    konst_1266_wire_constant <= "100";
    konst_1272_wire_constant <= "001";
    konst_1276_wire_constant <= "00000000000000000000000000000000";
    konst_1279_wire_constant <= "010";
    konst_1283_wire_constant <= "00000000000000000000000000000000";
    konst_1287_wire_constant <= "011";
    konst_1291_wire_constant <= "00000000000000000000000000000000";
    konst_1294_wire_constant <= "100";
    konst_1298_wire_constant <= "00000000000000000000000000000000";
    konst_1305_wire_constant <= "001";
    konst_1308_wire_constant <= "0";
    konst_1311_wire_constant <= "010";
    konst_1314_wire_constant <= "0";
    konst_1318_wire_constant <= "011";
    konst_1321_wire_constant <= "0";
    konst_1324_wire_constant <= "100";
    konst_1327_wire_constant <= "0";
    konst_1346_wire_constant <= "1";
    type_cast_1106_wire_constant <= "0";
    phi_stmt_1045: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_8_1047_wire_constant & next_down_counter_1237_1048_buffered;
      req <= phi_stmt_1045_req_0 & phi_stmt_1045_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1045",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1045_ack_0,
          idata => idata,
          odata => down_counter_1045,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1045
    phi_stmt_1049: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1051_wire_constant & RPIPE_noblock_obuf_1_1_1053_wire;
      req <= phi_stmt_1049_req_0 & phi_stmt_1049_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1049",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1049_ack_0,
          idata => idata,
          odata => pkt_1_e_word_1049,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1049
    phi_stmt_1054: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1056_wire_constant & RPIPE_noblock_obuf_2_1_1058_wire;
      req <= phi_stmt_1054_req_0 & phi_stmt_1054_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1054",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1054_ack_0,
          idata => idata,
          odata => pkt_2_e_word_1054,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1054
    phi_stmt_1059: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1061_wire_constant & RPIPE_noblock_obuf_3_1_1063_wire;
      req <= phi_stmt_1059_req_0 & phi_stmt_1059_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1059",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1059_ack_0,
          idata => idata,
          odata => pkt_3_e_word_1059,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1059
    phi_stmt_1064: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1066_wire_constant & RPIPE_noblock_obuf_4_1_1068_wire;
      req <= phi_stmt_1064_req_0 & phi_stmt_1064_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1064",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1064_ack_0,
          idata => idata,
          odata => pkt_4_e_word_1064,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1064
    phi_stmt_1069: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_3_1071_wire_constant & next_active_packet_1179_1072_buffered;
      req <= phi_stmt_1069_req_0 & phi_stmt_1069_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1069",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1069_ack_0,
          idata => idata,
          odata => active_packet_1069,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1069
    phi_stmt_1073: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_8_1075_wire_constant & next_active_packet_length_1224_1076_buffered;
      req <= phi_stmt_1073_req_0 & phi_stmt_1073_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1073",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1073_ack_0,
          idata => idata,
          odata => active_packet_length_1073,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1073
    phi_stmt_1077: Block -- phi operator 
      signal idata: std_logic_vector(3 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_2_1079_wire_constant & next_priority_index_1179_1080_buffered;
      req <= phi_stmt_1077_req_0 & phi_stmt_1077_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1077",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 2) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1077_ack_0,
          idata => idata,
          odata => priority_index_1077,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1077
    -- flow-through select operator MUX_1086_inst
    MUX_1086_wire <= konst_1084_wire_constant when (read_from_1_1245(0) /=  '0') else konst_1085_wire_constant;
    -- flow-through select operator MUX_1090_inst
    MUX_1090_wire <= konst_1088_wire_constant when (read_from_2_1253(0) /=  '0') else konst_1089_wire_constant;
    -- flow-through select operator MUX_1095_inst
    MUX_1095_wire <= konst_1093_wire_constant when (read_from_3_1261(0) /=  '0') else konst_1094_wire_constant;
    -- flow-through select operator MUX_1099_inst
    MUX_1099_wire <= konst_1097_wire_constant when (read_from_4_1269(0) /=  '0') else konst_1098_wire_constant;
    -- flow-through select operator MUX_1147_inst
    MUX_1147_wire <= p1_valid_1113 when (EQ_u3_u1_1144_wire(0) /=  '0') else konst_1146_wire_constant;
    -- flow-through select operator MUX_1153_inst
    MUX_1153_wire <= p2_valid_1118 when (EQ_u3_u1_1150_wire(0) /=  '0') else konst_1152_wire_constant;
    -- flow-through select operator MUX_1160_inst
    MUX_1160_wire <= p3_valid_1123 when (EQ_u3_u1_1157_wire(0) /=  '0') else konst_1159_wire_constant;
    -- flow-through select operator MUX_1166_inst
    MUX_1166_wire <= p4_valid_1128 when (EQ_u3_u1_1163_wire(0) /=  '0') else konst_1165_wire_constant;
    -- flow-through select operator MUX_1197_inst
    MUX_1197_wire <= slice_1195_wire when (EQ_u3_u1_1193_wire(0) /=  '0') else konst_1196_wire_constant;
    -- flow-through select operator MUX_1204_inst
    MUX_1204_wire <= slice_1202_wire when (EQ_u3_u1_1200_wire(0) /=  '0') else konst_1203_wire_constant;
    -- flow-through select operator MUX_1212_inst
    MUX_1212_wire <= slice_1210_wire when (EQ_u3_u1_1208_wire(0) /=  '0') else konst_1211_wire_constant;
    -- flow-through select operator MUX_1219_inst
    MUX_1219_wire <= slice_1217_wire when (EQ_u3_u1_1215_wire(0) /=  '0') else konst_1218_wire_constant;
    -- flow-through select operator MUX_1223_inst
    next_active_packet_length_1224 <= OR_u8_u8_1221_wire when (started_new_packet_1188(0) /=  '0') else active_packet_length_1073;
    -- flow-through select operator MUX_1235_inst
    MUX_1235_wire <= SUB_u8_u8_1233_wire when (valid_active_pkt_word_read_1169(0) /=  '0') else down_counter_1045;
    -- flow-through select operator MUX_1236_inst
    next_down_counter_1237 <= SUB_u8_u8_1229_wire when (started_new_packet_1188(0) /=  '0') else MUX_1235_wire;
    -- flow-through select operator MUX_1277_inst
    MUX_1277_wire <= slice_1275_wire when (EQ_u3_u1_1273_wire(0) /=  '0') else konst_1276_wire_constant;
    -- flow-through select operator MUX_1284_inst
    MUX_1284_wire <= slice_1282_wire when (EQ_u3_u1_1280_wire(0) /=  '0') else konst_1283_wire_constant;
    -- flow-through select operator MUX_1292_inst
    MUX_1292_wire <= slice_1290_wire when (EQ_u3_u1_1288_wire(0) /=  '0') else konst_1291_wire_constant;
    -- flow-through select operator MUX_1299_inst
    MUX_1299_wire <= slice_1297_wire when (EQ_u3_u1_1295_wire(0) /=  '0') else konst_1298_wire_constant;
    -- flow-through select operator MUX_1309_inst
    MUX_1309_wire <= p1_valid_1113 when (EQ_u3_u1_1306_wire(0) /=  '0') else konst_1308_wire_constant;
    -- flow-through select operator MUX_1315_inst
    MUX_1315_wire <= p2_valid_1118 when (EQ_u3_u1_1312_wire(0) /=  '0') else konst_1314_wire_constant;
    -- flow-through select operator MUX_1322_inst
    MUX_1322_wire <= p3_valid_1123 when (EQ_u3_u1_1319_wire(0) /=  '0') else konst_1321_wire_constant;
    -- flow-through select operator MUX_1328_inst
    MUX_1328_wire <= p4_valid_1128 when (EQ_u3_u1_1325_wire(0) /=  '0') else konst_1327_wire_constant;
    -- flow-through slice operator slice_1195_inst
    slice_1195_wire <= pkt_1_e_word_1049(15 downto 8);
    -- flow-through slice operator slice_1202_inst
    slice_1202_wire <= pkt_2_e_word_1054(15 downto 8);
    -- flow-through slice operator slice_1210_inst
    slice_1210_wire <= pkt_3_e_word_1059(15 downto 8);
    -- flow-through slice operator slice_1217_inst
    slice_1217_wire <= pkt_4_e_word_1064(15 downto 8);
    -- flow-through slice operator slice_1275_inst
    slice_1275_wire <= pkt_1_e_word_1049(31 downto 0);
    -- flow-through slice operator slice_1282_inst
    slice_1282_wire <= pkt_2_e_word_1054(31 downto 0);
    -- flow-through slice operator slice_1290_inst
    slice_1290_wire <= pkt_3_e_word_1059(31 downto 0);
    -- flow-through slice operator slice_1297_inst
    slice_1297_wire <= pkt_4_e_word_1064(31 downto 0);
    next_active_packet_1179_1072_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_active_packet_1179_1072_buf_req_0;
      next_active_packet_1179_1072_buf_ack_0<= wack(0);
      rreq(0) <= next_active_packet_1179_1072_buf_req_1;
      next_active_packet_1179_1072_buf_ack_1<= rack(0);
      next_active_packet_1179_1072_buf : InterlockBuffer generic map ( -- 
        name => "next_active_packet_1179_1072_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_active_packet_1179,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_active_packet_1179_1072_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_active_packet_length_1224_1076_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_active_packet_length_1224_1076_buf_req_0;
      next_active_packet_length_1224_1076_buf_ack_0<= wack(0);
      rreq(0) <= next_active_packet_length_1224_1076_buf_req_1;
      next_active_packet_length_1224_1076_buf_ack_1<= rack(0);
      next_active_packet_length_1224_1076_buf : InterlockBuffer generic map ( -- 
        name => "next_active_packet_length_1224_1076_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_active_packet_length_1224,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_active_packet_length_1224_1076_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_down_counter_1237_1048_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_down_counter_1237_1048_buf_req_0;
      next_down_counter_1237_1048_buf_ack_0<= wack(0);
      rreq(0) <= next_down_counter_1237_1048_buf_req_1;
      next_down_counter_1237_1048_buf_ack_1<= rack(0);
      next_down_counter_1237_1048_buf : InterlockBuffer generic map ( -- 
        name => "next_down_counter_1237_1048_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_down_counter_1237,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_down_counter_1237_1048_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_priority_index_1179_1080_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_priority_index_1179_1080_buf_req_0;
      next_priority_index_1179_1080_buf_ack_0<= wack(0);
      rreq(0) <= next_priority_index_1179_1080_buf_req_1;
      next_priority_index_1179_1080_buf_ack_1<= rack(0);
      next_priority_index_1179_1080_buf : InterlockBuffer generic map ( -- 
        name => "next_priority_index_1179_1080_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 2,
        out_data_width => 2,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_priority_index_1179,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_priority_index_1179_1080_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1043_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1346_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1043_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1043_branch_req_0,
          ack0 => do_while_stmt_1043_branch_ack_0,
          ack1 => do_while_stmt_1043_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- flow through binary operator AND_u1_u1_1187_inst
    started_new_packet_1188 <= (NEQ_u3_u1_1183_wire and EQ_u8_u1_1186_wire);
    -- flow through binary operator BITSEL_u33_u1_1112_inst
    process(pkt_1_e_word_1049) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_1_e_word_1049, konst_1111_wire_constant, tmp_var);
      p1_valid_1113 <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u33_u1_1117_inst
    process(pkt_2_e_word_1054) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_2_e_word_1054, konst_1116_wire_constant, tmp_var);
      p2_valid_1118 <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u33_u1_1122_inst
    process(pkt_3_e_word_1059) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_3_e_word_1059, konst_1121_wire_constant, tmp_var);
      p3_valid_1123 <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u33_u1_1127_inst
    process(pkt_4_e_word_1064) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_4_e_word_1064, konst_1126_wire_constant, tmp_var);
      p4_valid_1128 <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1144_inst
    process(active_packet_1069) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1069, konst_1143_wire_constant, tmp_var);
      EQ_u3_u1_1144_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1150_inst
    process(active_packet_1069) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1069, konst_1149_wire_constant, tmp_var);
      EQ_u3_u1_1150_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1157_inst
    process(active_packet_1069) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1069, konst_1156_wire_constant, tmp_var);
      EQ_u3_u1_1157_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1163_inst
    process(active_packet_1069) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1069, konst_1162_wire_constant, tmp_var);
      EQ_u3_u1_1163_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1193_inst
    process(next_active_packet_1179) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1179, konst_1192_wire_constant, tmp_var);
      EQ_u3_u1_1193_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1200_inst
    process(next_active_packet_1179) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1179, konst_1199_wire_constant, tmp_var);
      EQ_u3_u1_1200_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1208_inst
    process(next_active_packet_1179) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1179, konst_1207_wire_constant, tmp_var);
      EQ_u3_u1_1208_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1215_inst
    process(next_active_packet_1179) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1179, konst_1214_wire_constant, tmp_var);
      EQ_u3_u1_1215_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1243_inst
    process(next_active_packet_1179) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1179, konst_1242_wire_constant, tmp_var);
      EQ_u3_u1_1243_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1251_inst
    process(next_active_packet_1179) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1179, konst_1250_wire_constant, tmp_var);
      EQ_u3_u1_1251_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1259_inst
    process(next_active_packet_1179) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1179, konst_1258_wire_constant, tmp_var);
      EQ_u3_u1_1259_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1267_inst
    process(next_active_packet_1179) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1179, konst_1266_wire_constant, tmp_var);
      EQ_u3_u1_1267_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1273_inst
    process(next_active_packet_1179) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1179, konst_1272_wire_constant, tmp_var);
      EQ_u3_u1_1273_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1280_inst
    process(next_active_packet_1179) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1179, konst_1279_wire_constant, tmp_var);
      EQ_u3_u1_1280_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1288_inst
    process(next_active_packet_1179) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1179, konst_1287_wire_constant, tmp_var);
      EQ_u3_u1_1288_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1295_inst
    process(next_active_packet_1179) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1179, konst_1294_wire_constant, tmp_var);
      EQ_u3_u1_1295_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1306_inst
    process(next_active_packet_1179) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1179, konst_1305_wire_constant, tmp_var);
      EQ_u3_u1_1306_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1312_inst
    process(next_active_packet_1179) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1179, konst_1311_wire_constant, tmp_var);
      EQ_u3_u1_1312_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1319_inst
    process(next_active_packet_1179) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1179, konst_1318_wire_constant, tmp_var);
      EQ_u3_u1_1319_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1325_inst
    process(next_active_packet_1179) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1179, konst_1324_wire_constant, tmp_var);
      EQ_u3_u1_1325_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u8_u1_1186_inst
    process(down_counter_1045) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(down_counter_1045, konst_1185_wire_constant, tmp_var);
      EQ_u8_u1_1186_wire <= tmp_var; --
    end process;
    -- flow through binary operator NEQ_u3_u1_1183_inst
    process(next_active_packet_1179) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(next_active_packet_1179, konst_1182_wire_constant, tmp_var);
      NEQ_u3_u1_1183_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1240_inst
    process(p1_valid_1113) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p1_valid_1113, tmp_var);
      NOT_u1_u1_1240_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1248_inst
    process(p2_valid_1118) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p2_valid_1118, tmp_var);
      NOT_u1_u1_1248_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1256_inst
    process(p3_valid_1123) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p3_valid_1123, tmp_var);
      NOT_u1_u1_1256_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1264_inst
    process(p4_valid_1128) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p4_valid_1128, tmp_var);
      NOT_u1_u1_1264_wire <= tmp_var; -- 
    end process;
    -- flow through binary operator OR_u1_u1_1154_inst
    OR_u1_u1_1154_wire <= (MUX_1147_wire or MUX_1153_wire);
    -- flow through binary operator OR_u1_u1_1167_inst
    OR_u1_u1_1167_wire <= (MUX_1160_wire or MUX_1166_wire);
    -- flow through binary operator OR_u1_u1_1168_inst
    valid_active_pkt_word_read_1169 <= (OR_u1_u1_1154_wire or OR_u1_u1_1167_wire);
    -- flow through binary operator OR_u1_u1_1244_inst
    read_from_1_1245 <= (NOT_u1_u1_1240_wire or EQ_u3_u1_1243_wire);
    -- flow through binary operator OR_u1_u1_1252_inst
    read_from_2_1253 <= (NOT_u1_u1_1248_wire or EQ_u3_u1_1251_wire);
    -- flow through binary operator OR_u1_u1_1260_inst
    read_from_3_1261 <= (NOT_u1_u1_1256_wire or EQ_u3_u1_1259_wire);
    -- flow through binary operator OR_u1_u1_1268_inst
    read_from_4_1269 <= (NOT_u1_u1_1264_wire or EQ_u3_u1_1267_wire);
    -- flow through binary operator OR_u1_u1_1316_inst
    OR_u1_u1_1316_wire <= (MUX_1309_wire or MUX_1315_wire);
    -- flow through binary operator OR_u1_u1_1329_inst
    OR_u1_u1_1329_wire <= (MUX_1322_wire or MUX_1328_wire);
    -- flow through binary operator OR_u1_u1_1330_inst
    send_flag_1331 <= (OR_u1_u1_1316_wire or OR_u1_u1_1329_wire);
    -- flow through binary operator OR_u32_u32_1285_inst
    OR_u32_u32_1285_wire <= (MUX_1277_wire or MUX_1284_wire);
    -- flow through binary operator OR_u32_u32_1300_inst
    OR_u32_u32_1300_wire <= (MUX_1292_wire or MUX_1299_wire);
    -- flow through binary operator OR_u32_u32_1301_inst
    data_to_out_1302 <= (OR_u32_u32_1285_wire or OR_u32_u32_1300_wire);
    -- flow through binary operator OR_u8_u8_1091_inst
    OR_u8_u8_1091_wire <= (MUX_1086_wire or MUX_1090_wire);
    -- flow through binary operator OR_u8_u8_1100_inst
    OR_u8_u8_1100_wire <= (MUX_1095_wire or MUX_1099_wire);
    -- flow through binary operator OR_u8_u8_1101_inst
    senderPort_1102 <= (OR_u8_u8_1091_wire or OR_u8_u8_1100_wire);
    -- flow through binary operator OR_u8_u8_1205_inst
    OR_u8_u8_1205_wire <= (MUX_1197_wire or MUX_1204_wire);
    -- flow through binary operator OR_u8_u8_1220_inst
    OR_u8_u8_1220_wire <= (MUX_1212_wire or MUX_1219_wire);
    -- flow through binary operator OR_u8_u8_1221_inst
    OR_u8_u8_1221_wire <= (OR_u8_u8_1205_wire or OR_u8_u8_1220_wire);
    -- flow through binary operator SUB_u8_u8_1229_inst
    SUB_u8_u8_1229_wire <= std_logic_vector(unsigned(next_active_packet_length_1224) - unsigned(konst_1228_wire_constant));
    -- flow through binary operator SUB_u8_u8_1233_inst
    SUB_u8_u8_1233_wire <= std_logic_vector(unsigned(down_counter_1045) - unsigned(konst_1232_wire_constant));
    -- shared inport operator group (0) : RPIPE_noblock_obuf_1_1_1053_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_1_1_1053_inst_req_0;
      RPIPE_noblock_obuf_1_1_1053_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_1_1_1053_inst_req_1;
      RPIPE_noblock_obuf_1_1_1053_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_1_1245(0);
      RPIPE_noblock_obuf_1_1_1053_wire <= data_out(32 downto 0);
      noblock_obuf_1_1_read_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_1_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_1_read_0: InputPortRevised -- 
        generic map ( name => "noblock_obuf_1_1_read_0", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_1_1_pipe_read_req(0),
          oack => noblock_obuf_1_1_pipe_read_ack(0),
          odata => noblock_obuf_1_1_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_noblock_obuf_2_1_1058_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_2_1_1058_inst_req_0;
      RPIPE_noblock_obuf_2_1_1058_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_2_1_1058_inst_req_1;
      RPIPE_noblock_obuf_2_1_1058_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_2_1253(0);
      RPIPE_noblock_obuf_2_1_1058_wire <= data_out(32 downto 0);
      noblock_obuf_2_1_read_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_1_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_1_read_1: InputPortRevised -- 
        generic map ( name => "noblock_obuf_2_1_read_1", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_2_1_pipe_read_req(0),
          oack => noblock_obuf_2_1_pipe_read_ack(0),
          odata => noblock_obuf_2_1_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_noblock_obuf_3_1_1063_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_3_1_1063_inst_req_0;
      RPIPE_noblock_obuf_3_1_1063_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_3_1_1063_inst_req_1;
      RPIPE_noblock_obuf_3_1_1063_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_3_1261(0);
      RPIPE_noblock_obuf_3_1_1063_wire <= data_out(32 downto 0);
      noblock_obuf_3_1_read_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_1_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_1_read_2: InputPortRevised -- 
        generic map ( name => "noblock_obuf_3_1_read_2", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_3_1_pipe_read_req(0),
          oack => noblock_obuf_3_1_pipe_read_ack(0),
          odata => noblock_obuf_3_1_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_noblock_obuf_4_1_1068_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_4_1_1068_inst_req_0;
      RPIPE_noblock_obuf_4_1_1068_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_4_1_1068_inst_req_1;
      RPIPE_noblock_obuf_4_1_1068_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_4_1269(0);
      RPIPE_noblock_obuf_4_1_1068_wire <= data_out(32 downto 0);
      noblock_obuf_4_1_read_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_1_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_1_read_3: InputPortRevised -- 
        generic map ( name => "noblock_obuf_4_1_read_3", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_4_1_pipe_read_req(0),
          oack => noblock_obuf_4_1_pipe_read_ack(0),
          odata => noblock_obuf_4_1_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_out_data_1_1333_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_out_data_1_1333_inst_req_0;
      WPIPE_out_data_1_1333_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_out_data_1_1333_inst_req_1;
      WPIPE_out_data_1_1333_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_flag_1331(0);
      data_in <= data_to_out_1302;
      out_data_1_write_0_gI: SplitGuardInterface generic map(name => "out_data_1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      out_data_1_write_0: OutputPortRevised -- 
        generic map ( name => "out_data_1", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => out_data_1_pipe_write_req(0),
          oack => out_data_1_pipe_write_ack(0),
          odata => out_data_1_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_1108_call 
    updateCounter_call_group_0: Block -- 
      signal data_in: std_logic_vector(16 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1108_call_req_0;
      call_stmt_1108_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1108_call_req_1;
      call_stmt_1108_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      updateCounter_call_group_0_gI: SplitGuardInterface generic map(name => "updateCounter_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= senderPort_1102 & konst_1104_wire_constant & type_cast_1106_wire_constant;
      continue_1108 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 17,
        owidth => 17,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => updateCounter_call_reqs(0),
          ackR => updateCounter_call_acks(0),
          dataR => updateCounter_call_data(16 downto 0),
          tagR => updateCounter_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => updateCounter_return_acks(0), -- cross-over
          ackL => updateCounter_return_reqs(0), -- cross-over
          dataL => updateCounter_return_data(0 downto 0),
          tagL => updateCounter_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    volatile_operator_prioritySelect_4206: prioritySelect_Volatile port map(down_counter => down_counter_1045, active_packet => active_packet_1069, priority_index => priority_index_1077, p1_valid => p1_valid_1113, p2_valid => p2_valid_1118, p3_valid => p3_valid_1123, p4_valid => p4_valid_1128, next_active_packet => next_active_packet_1179, next_priority_index => next_priority_index_1179); 
    -- 
  end Block; -- data_path
  -- 
end outputPort_1_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity outputPort_2_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    noblock_obuf_1_2_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_2_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_3_2_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_2_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_4_2_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_2_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_2_2_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_2_pipe_read_data : in   std_logic_vector(32 downto 0);
    out_data_2_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_data_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_data_2_pipe_write_data : out  std_logic_vector(31 downto 0);
    updateCounter_call_reqs : out  std_logic_vector(0 downto 0);
    updateCounter_call_acks : in   std_logic_vector(0 downto 0);
    updateCounter_call_data : out  std_logic_vector(16 downto 0);
    updateCounter_call_tag  :  out  std_logic_vector(0 downto 0);
    updateCounter_return_reqs : out  std_logic_vector(0 downto 0);
    updateCounter_return_acks : in   std_logic_vector(0 downto 0);
    updateCounter_return_data : in   std_logic_vector(0 downto 0);
    updateCounter_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity outputPort_2_Daemon;
architecture outputPort_2_Daemon_arch of outputPort_2_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal outputPort_2_Daemon_CP_2845_start: Boolean;
  signal outputPort_2_Daemon_CP_2845_symbol: Boolean;
  -- volatile/operator module components. 
  component updateCounter is -- 
    generic (tag_length : integer); 
    port ( -- 
      input_port : in  std_logic_vector(7 downto 0);
      output_port : in  std_logic_vector(7 downto 0);
      up : in  std_logic_vector(0 downto 0);
      continue : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(3 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(1 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(1 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component prioritySelect_Volatile is -- 
    port ( -- 
      down_counter : in  std_logic_vector(7 downto 0);
      active_packet : in  std_logic_vector(2 downto 0);
      priority_index : in  std_logic_vector(1 downto 0);
      p1_valid : in  std_logic_vector(0 downto 0);
      p2_valid : in  std_logic_vector(0 downto 0);
      p3_valid : in  std_logic_vector(0 downto 0);
      p4_valid : in  std_logic_vector(0 downto 0);
      next_active_packet : out  std_logic_vector(2 downto 0);
      next_priority_index : out  std_logic_vector(1 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal next_down_counter_1545_1356_buf_ack_1 : boolean;
  signal next_down_counter_1545_1356_buf_req_0 : boolean;
  signal next_down_counter_1545_1356_buf_ack_0 : boolean;
  signal call_stmt_1416_call_req_1 : boolean;
  signal phi_stmt_1353_req_0 : boolean;
  signal phi_stmt_1353_req_1 : boolean;
  signal call_stmt_1416_call_ack_1 : boolean;
  signal do_while_stmt_1351_branch_req_0 : boolean;
  signal phi_stmt_1353_ack_0 : boolean;
  signal next_down_counter_1545_1356_buf_req_1 : boolean;
  signal WPIPE_out_data_2_1641_inst_req_0 : boolean;
  signal WPIPE_out_data_2_1641_inst_ack_0 : boolean;
  signal WPIPE_out_data_2_1641_inst_req_1 : boolean;
  signal WPIPE_out_data_2_1641_inst_ack_1 : boolean;
  signal do_while_stmt_1351_branch_ack_0 : boolean;
  signal do_while_stmt_1351_branch_ack_1 : boolean;
  signal phi_stmt_1385_ack_0 : boolean;
  signal phi_stmt_1385_req_0 : boolean;
  signal phi_stmt_1357_req_1 : boolean;
  signal phi_stmt_1357_req_0 : boolean;
  signal call_stmt_1416_call_ack_0 : boolean;
  signal call_stmt_1416_call_req_0 : boolean;
  signal phi_stmt_1357_ack_0 : boolean;
  signal phi_stmt_1367_ack_0 : boolean;
  signal phi_stmt_1385_req_1 : boolean;
  signal next_priority_index_1487_1388_buf_ack_1 : boolean;
  signal next_priority_index_1487_1388_buf_req_1 : boolean;
  signal next_priority_index_1487_1388_buf_ack_0 : boolean;
  signal next_priority_index_1487_1388_buf_req_0 : boolean;
  signal RPIPE_noblock_obuf_1_2_1361_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_1_2_1361_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_1_2_1361_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_1_2_1361_inst_ack_1 : boolean;
  signal phi_stmt_1362_req_1 : boolean;
  signal phi_stmt_1362_req_0 : boolean;
  signal phi_stmt_1362_ack_0 : boolean;
  signal RPIPE_noblock_obuf_2_2_1366_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_2_2_1366_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_2_2_1366_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_2_2_1366_inst_ack_1 : boolean;
  signal phi_stmt_1367_req_1 : boolean;
  signal phi_stmt_1367_req_0 : boolean;
  signal RPIPE_noblock_obuf_3_2_1371_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_3_2_1371_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_3_2_1371_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_3_2_1371_inst_ack_1 : boolean;
  signal phi_stmt_1372_req_1 : boolean;
  signal phi_stmt_1372_req_0 : boolean;
  signal phi_stmt_1372_ack_0 : boolean;
  signal RPIPE_noblock_obuf_4_2_1376_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_4_2_1376_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_4_2_1376_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_4_2_1376_inst_ack_1 : boolean;
  signal phi_stmt_1377_req_1 : boolean;
  signal phi_stmt_1377_req_0 : boolean;
  signal phi_stmt_1377_ack_0 : boolean;
  signal next_active_packet_1487_1380_buf_req_0 : boolean;
  signal next_active_packet_1487_1380_buf_ack_0 : boolean;
  signal next_active_packet_1487_1380_buf_req_1 : boolean;
  signal next_active_packet_1487_1380_buf_ack_1 : boolean;
  signal phi_stmt_1381_req_1 : boolean;
  signal phi_stmt_1381_req_0 : boolean;
  signal phi_stmt_1381_ack_0 : boolean;
  signal next_active_packet_length_1532_1384_buf_req_0 : boolean;
  signal next_active_packet_length_1532_1384_buf_ack_0 : boolean;
  signal next_active_packet_length_1532_1384_buf_req_1 : boolean;
  signal next_active_packet_length_1532_1384_buf_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "outputPort_2_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  outputPort_2_Daemon_CP_2845_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "outputPort_2_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_2_Daemon_CP_2845_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= outputPort_2_Daemon_CP_2845_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_2_Daemon_CP_2845_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  outputPort_2_Daemon_CP_2845: Block -- control-path 
    signal outputPort_2_Daemon_CP_2845_elements: BooleanArray(185 downto 0);
    -- 
  begin -- 
    outputPort_2_Daemon_CP_2845_elements(0) <= outputPort_2_Daemon_CP_2845_start;
    outputPort_2_Daemon_CP_2845_symbol <= outputPort_2_Daemon_CP_2845_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1350/branch_block_stmt_1350__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1350/$entry
      -- CP-element group 0: 	 branch_block_stmt_1350/do_while_stmt_1351__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	185 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1350/branch_block_stmt_1350__exit__
      -- CP-element group 1: 	 branch_block_stmt_1350/$exit
      -- CP-element group 1: 	 branch_block_stmt_1350/do_while_stmt_1351__exit__
      -- 
    outputPort_2_Daemon_CP_2845_elements(1) <= outputPort_2_Daemon_CP_2845_elements(185);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1350/do_while_stmt_1351/$entry
      -- CP-element group 2: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351__entry__
      -- 
    outputPort_2_Daemon_CP_2845_elements(2) <= outputPort_2_Daemon_CP_2845_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	185 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351__exit__
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1350/do_while_stmt_1351/loop_back
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	184 
    -- CP-element group 5: 	183 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1350/do_while_stmt_1351/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1350/do_while_stmt_1351/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1350/do_while_stmt_1351/loop_taken/$entry
      -- 
    outputPort_2_Daemon_CP_2845_elements(5) <= outputPort_2_Daemon_CP_2845_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	182 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1350/do_while_stmt_1351/loop_body_done
      -- 
    outputPort_2_Daemon_CP_2845_elements(6) <= outputPort_2_Daemon_CP_2845_elements(182);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	143 
    -- CP-element group 7: 	161 
    -- CP-element group 7: 	22 
    -- CP-element group 7: 	41 
    -- CP-element group 7: 	62 
    -- CP-element group 7: 	83 
    -- CP-element group 7: 	104 
    -- CP-element group 7: 	125 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/back_edge_to_loop_body
      -- 
    outputPort_2_Daemon_CP_2845_elements(7) <= outputPort_2_Daemon_CP_2845_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	163 
    -- CP-element group 8: 	145 
    -- CP-element group 8: 	24 
    -- CP-element group 8: 	43 
    -- CP-element group 8: 	64 
    -- CP-element group 8: 	85 
    -- CP-element group 8: 	106 
    -- CP-element group 8: 	127 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/first_time_through_loop_body
      -- 
    outputPort_2_Daemon_CP_2845_elements(8) <= outputPort_2_Daemon_CP_2845_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	157 
    -- CP-element group 9: 	181 
    -- CP-element group 9: 	156 
    -- CP-element group 9: 	139 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	17 
    -- CP-element group 9: 	35 
    -- CP-element group 9: 	36 
    -- CP-element group 9: 	56 
    -- CP-element group 9: 	57 
    -- CP-element group 9: 	77 
    -- CP-element group 9: 	78 
    -- CP-element group 9: 	98 
    -- CP-element group 9: 	99 
    -- CP-element group 9: 	119 
    -- CP-element group 9: 	120 
    -- CP-element group 9: 	138 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/loop_body_start
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	181 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/condition_evaluated
      -- 
    condition_evaluated_2869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(10), ack => do_while_stmt_1351_branch_req_0); -- 
    outputPort_2_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(181) & outputPort_2_Daemon_CP_2845_elements(15);
      gj_outputPort_2_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	156 
    -- CP-element group 11: 	16 
    -- CP-element group 11: 	35 
    -- CP-element group 11: 	56 
    -- CP-element group 11: 	77 
    -- CP-element group 11: 	98 
    -- CP-element group 11: 	119 
    -- CP-element group 11: 	138 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	158 
    -- CP-element group 11: 	18 
    -- CP-element group 11: 	37 
    -- CP-element group 11: 	58 
    -- CP-element group 11: 	79 
    -- CP-element group 11: 	100 
    -- CP-element group 11: 	121 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1381_sample_start__ps
      -- 
    outputPort_2_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 1);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(156) & outputPort_2_Daemon_CP_2845_elements(16) & outputPort_2_Daemon_CP_2845_elements(35) & outputPort_2_Daemon_CP_2845_elements(56) & outputPort_2_Daemon_CP_2845_elements(77) & outputPort_2_Daemon_CP_2845_elements(98) & outputPort_2_Daemon_CP_2845_elements(119) & outputPort_2_Daemon_CP_2845_elements(138) & outputPort_2_Daemon_CP_2845_elements(15);
      gj_outputPort_2_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	140 
    -- CP-element group 12: 	159 
    -- CP-element group 12: 	19 
    -- CP-element group 12: 	38 
    -- CP-element group 12: 	59 
    -- CP-element group 12: 	80 
    -- CP-element group 12: 	101 
    -- CP-element group 12: 	122 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	182 
    -- CP-element group 12: 	13 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	156 
    -- CP-element group 12: 	16 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	56 
    -- CP-element group 12: 	77 
    -- CP-element group 12: 	98 
    -- CP-element group 12: 	119 
    -- CP-element group 12: 	138 
    -- CP-element group 12:  members (9) 
      -- CP-element group 12: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1353_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1357_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1362_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1367_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1372_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1377_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1381_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1385_sample_completed_
      -- 
    outputPort_2_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(140) & outputPort_2_Daemon_CP_2845_elements(159) & outputPort_2_Daemon_CP_2845_elements(19) & outputPort_2_Daemon_CP_2845_elements(38) & outputPort_2_Daemon_CP_2845_elements(59) & outputPort_2_Daemon_CP_2845_elements(80) & outputPort_2_Daemon_CP_2845_elements(101) & outputPort_2_Daemon_CP_2845_elements(122);
      gj_outputPort_2_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	182 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/aggregated_phi_sample_ack_d
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(13) is a control-delay.
    cp_element_13_delay: control_delay_element  generic map(name => " 13_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_2845_elements(12), ack => outputPort_2_Daemon_CP_2845_elements(13), clk => clk, reset =>reset);
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	157 
    -- CP-element group 14: 	139 
    -- CP-element group 14: 	17 
    -- CP-element group 14: 	36 
    -- CP-element group 14: 	57 
    -- CP-element group 14: 	78 
    -- CP-element group 14: 	99 
    -- CP-element group 14: 	120 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	141 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	39 
    -- CP-element group 14: 	60 
    -- CP-element group 14: 	81 
    -- CP-element group 14: 	102 
    -- CP-element group 14: 	123 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/aggregated_phi_update_req
      -- CP-element group 14: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1385_update_start__ps
      -- 
    outputPort_2_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(157) & outputPort_2_Daemon_CP_2845_elements(139) & outputPort_2_Daemon_CP_2845_elements(17) & outputPort_2_Daemon_CP_2845_elements(36) & outputPort_2_Daemon_CP_2845_elements(57) & outputPort_2_Daemon_CP_2845_elements(78) & outputPort_2_Daemon_CP_2845_elements(99) & outputPort_2_Daemon_CP_2845_elements(120);
      gj_outputPort_2_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	160 
    -- CP-element group 15: 	142 
    -- CP-element group 15: 	21 
    -- CP-element group 15: 	40 
    -- CP-element group 15: 	61 
    -- CP-element group 15: 	82 
    -- CP-element group 15: 	103 
    -- CP-element group 15: 	124 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/aggregated_phi_update_ack
      -- 
    outputPort_2_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 7);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(160) & outputPort_2_Daemon_CP_2845_elements(142) & outputPort_2_Daemon_CP_2845_elements(21) & outputPort_2_Daemon_CP_2845_elements(40) & outputPort_2_Daemon_CP_2845_elements(61) & outputPort_2_Daemon_CP_2845_elements(82) & outputPort_2_Daemon_CP_2845_elements(103) & outputPort_2_Daemon_CP_2845_elements(124);
      gj_outputPort_2_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	11 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1353_sample_start_
      -- 
    outputPort_2_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(9) & outputPort_2_Daemon_CP_2845_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	9 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	176 
    -- CP-element group 17: 	179 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	14 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1353_update_start_
      -- 
    outputPort_2_Daemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(9) & outputPort_2_Daemon_CP_2845_elements(176) & outputPort_2_Daemon_CP_2845_elements(179);
      gj_outputPort_2_Daemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	11 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1353_sample_start__ps
      -- 
    outputPort_2_Daemon_CP_2845_elements(18) <= outputPort_2_Daemon_CP_2845_elements(11);
    -- CP-element group 19:  join  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	12 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1353_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(19) is bound as output of CP function.
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	14 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1353_update_start__ps
      -- 
    outputPort_2_Daemon_CP_2845_elements(20) <= outputPort_2_Daemon_CP_2845_elements(14);
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	174 
    -- CP-element group 21: 	178 
    -- CP-element group 21: 	15 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1353_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1353_update_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(21) is bound as output of CP function.
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	7 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1353_loopback_trigger
      -- 
    outputPort_2_Daemon_CP_2845_elements(22) <= outputPort_2_Daemon_CP_2845_elements(7);
    -- CP-element group 23:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1353_loopback_sample_req_ps
      -- CP-element group 23: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1353_loopback_sample_req
      -- 
    phi_stmt_1353_loopback_sample_req_2885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1353_loopback_sample_req_2885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(23), ack => phi_stmt_1353_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(23) is bound as output of CP function.
    -- CP-element group 24:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	8 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1353_entry_trigger
      -- 
    outputPort_2_Daemon_CP_2845_elements(24) <= outputPort_2_Daemon_CP_2845_elements(8);
    -- CP-element group 25:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1353_entry_sample_req
      -- CP-element group 25: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1353_entry_sample_req_ps
      -- 
    phi_stmt_1353_entry_sample_req_2888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1353_entry_sample_req_2888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(25), ack => phi_stmt_1353_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1353_phi_mux_ack_ps
      -- CP-element group 26: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1353_phi_mux_ack
      -- 
    phi_stmt_1353_phi_mux_ack_2891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1353_ack_0, ack => outputPort_2_Daemon_CP_2845_elements(26)); -- 
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_8_1355_sample_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_8_1355_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_8_1355_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_8_1355_sample_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_8_1355_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_8_1355_update_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	30 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_8_1355_update_completed__ps
      -- 
    outputPort_2_Daemon_CP_2845_elements(29) <= outputPort_2_Daemon_CP_2845_elements(30);
    -- CP-element group 30:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	29 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_8_1355_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(30) is a control-delay.
    cp_element_30_delay: control_delay_element  generic map(name => " 30_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_2845_elements(28), ack => outputPort_2_Daemon_CP_2845_elements(30), clk => clk, reset =>reset);
    -- CP-element group 31:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_down_counter_1356_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_down_counter_1356_Sample/req
      -- CP-element group 31: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_down_counter_1356_sample_start__ps
      -- CP-element group 31: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_down_counter_1356_sample_start_
      -- 
    req_2912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(31), ack => next_down_counter_1545_1356_buf_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_down_counter_1356_update_start__ps
      -- CP-element group 32: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_down_counter_1356_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_down_counter_1356_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_down_counter_1356_Update/req
      -- 
    req_2917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(32), ack => next_down_counter_1545_1356_buf_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_down_counter_1356_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_down_counter_1356_Sample/ack
      -- CP-element group 33: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_down_counter_1356_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_down_counter_1356_sample_completed__ps
      -- 
    ack_2913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_1545_1356_buf_ack_0, ack => outputPort_2_Daemon_CP_2845_elements(33)); -- 
    -- CP-element group 34:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_down_counter_1356_Update/ack
      -- CP-element group 34: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_down_counter_1356_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_down_counter_1356_update_completed__ps
      -- CP-element group 34: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_down_counter_1356_update_completed_
      -- 
    ack_2918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_1545_1356_buf_ack_1, ack => outputPort_2_Daemon_CP_2845_elements(34)); -- 
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	12 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	11 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1357_sample_start_
      -- 
    outputPort_2_Daemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(9) & outputPort_2_Daemon_CP_2845_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	9 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	176 
    -- CP-element group 36: 	179 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	14 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1357_update_start_
      -- 
    outputPort_2_Daemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(9) & outputPort_2_Daemon_CP_2845_elements(176) & outputPort_2_Daemon_CP_2845_elements(179);
      gj_outputPort_2_Daemon_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	11 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1357_sample_start__ps
      -- 
    outputPort_2_Daemon_CP_2845_elements(37) <= outputPort_2_Daemon_CP_2845_elements(11);
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	12 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1357_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(38) is bound as output of CP function.
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	14 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1357_update_start__ps
      -- 
    outputPort_2_Daemon_CP_2845_elements(39) <= outputPort_2_Daemon_CP_2845_elements(14);
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	174 
    -- CP-element group 40: 	178 
    -- CP-element group 40: 	15 
    -- CP-element group 40:  members (2) 
      -- CP-element group 40: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1357_update_completed__ps
      -- CP-element group 40: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1357_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(40) is bound as output of CP function.
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	7 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1357_loopback_trigger
      -- 
    outputPort_2_Daemon_CP_2845_elements(41) <= outputPort_2_Daemon_CP_2845_elements(7);
    -- CP-element group 42:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1357_loopback_sample_req
      -- CP-element group 42: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1357_loopback_sample_req_ps
      -- 
    phi_stmt_1357_loopback_sample_req_2929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1357_loopback_sample_req_2929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(42), ack => phi_stmt_1357_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(42) is bound as output of CP function.
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	8 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1357_entry_trigger
      -- 
    outputPort_2_Daemon_CP_2845_elements(43) <= outputPort_2_Daemon_CP_2845_elements(8);
    -- CP-element group 44:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1357_entry_sample_req
      -- CP-element group 44: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1357_entry_sample_req_ps
      -- 
    phi_stmt_1357_entry_sample_req_2932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1357_entry_sample_req_2932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(44), ack => phi_stmt_1357_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(44) is bound as output of CP function.
    -- CP-element group 45:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1357_phi_mux_ack
      -- CP-element group 45: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1357_phi_mux_ack_ps
      -- 
    phi_stmt_1357_phi_mux_ack_2935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1357_ack_0, ack => outputPort_2_Daemon_CP_2845_elements(45)); -- 
    -- CP-element group 46:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (4) 
      -- CP-element group 46: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1359_sample_start__ps
      -- CP-element group 46: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1359_sample_completed__ps
      -- CP-element group 46: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1359_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1359_sample_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1359_update_start__ps
      -- CP-element group 47: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1359_update_start_
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	49 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1359_update_completed__ps
      -- 
    outputPort_2_Daemon_CP_2845_elements(48) <= outputPort_2_Daemon_CP_2845_elements(49);
    -- CP-element group 49:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	48 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1359_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(49) is a control-delay.
    cp_element_49_delay: control_delay_element  generic map(name => " 49_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_2845_elements(47), ack => outputPort_2_Daemon_CP_2845_elements(49), clk => clk, reset =>reset);
    -- CP-element group 50:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_1_2_1361_sample_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_1_2_1361_update_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(51) is bound as output of CP function.
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	55 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_1_2_1361_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_1_2_1361_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_1_2_1361_Sample/rr
      -- 
    rr_2956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(52), ack => RPIPE_noblock_obuf_1_2_1361_inst_req_0); -- 
    outputPort_2_Daemon_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(50) & outputPort_2_Daemon_CP_2845_elements(55);
      gj_outputPort_2_Daemon_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: 	54 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_1_2_1361_update_start_
      -- CP-element group 53: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_1_2_1361_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_1_2_1361_Update/cr
      -- 
    cr_2961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(53), ack => RPIPE_noblock_obuf_1_2_1361_inst_req_1); -- 
    outputPort_2_Daemon_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(51) & outputPort_2_Daemon_CP_2845_elements(54);
      gj_outputPort_2_Daemon_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	53 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_1_2_1361_sample_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_1_2_1361_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_1_2_1361_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_1_2_1361_Sample/ra
      -- 
    ra_2957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_2_1361_inst_ack_0, ack => outputPort_2_Daemon_CP_2845_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: marked-successors 
    -- CP-element group 55: 	52 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_1_2_1361_update_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_1_2_1361_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_1_2_1361_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_1_2_1361_Update/ca
      -- 
    ca_2962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_2_1361_inst_ack_1, ack => outputPort_2_Daemon_CP_2845_elements(55)); -- 
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	9 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	12 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	11 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1362_sample_start_
      -- 
    outputPort_2_Daemon_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(9) & outputPort_2_Daemon_CP_2845_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  join  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	9 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	176 
    -- CP-element group 57: 	179 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	14 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1362_update_start_
      -- 
    outputPort_2_Daemon_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(9) & outputPort_2_Daemon_CP_2845_elements(176) & outputPort_2_Daemon_CP_2845_elements(179);
      gj_outputPort_2_Daemon_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	11 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1362_sample_start__ps
      -- 
    outputPort_2_Daemon_CP_2845_elements(58) <= outputPort_2_Daemon_CP_2845_elements(11);
    -- CP-element group 59:  join  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	12 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1362_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(59) is bound as output of CP function.
    -- CP-element group 60:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	14 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1362_update_start__ps
      -- 
    outputPort_2_Daemon_CP_2845_elements(60) <= outputPort_2_Daemon_CP_2845_elements(14);
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	174 
    -- CP-element group 61: 	178 
    -- CP-element group 61: 	15 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1362_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1362_update_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(61) is bound as output of CP function.
    -- CP-element group 62:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	7 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1362_loopback_trigger
      -- 
    outputPort_2_Daemon_CP_2845_elements(62) <= outputPort_2_Daemon_CP_2845_elements(7);
    -- CP-element group 63:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1362_loopback_sample_req
      -- CP-element group 63: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1362_loopback_sample_req_ps
      -- 
    phi_stmt_1362_loopback_sample_req_2973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1362_loopback_sample_req_2973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(63), ack => phi_stmt_1362_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(63) is bound as output of CP function.
    -- CP-element group 64:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	8 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1362_entry_trigger
      -- 
    outputPort_2_Daemon_CP_2845_elements(64) <= outputPort_2_Daemon_CP_2845_elements(8);
    -- CP-element group 65:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1362_entry_sample_req
      -- CP-element group 65: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1362_entry_sample_req_ps
      -- 
    phi_stmt_1362_entry_sample_req_2976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1362_entry_sample_req_2976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(65), ack => phi_stmt_1362_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(65) is bound as output of CP function.
    -- CP-element group 66:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1362_phi_mux_ack
      -- CP-element group 66: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1362_phi_mux_ack_ps
      -- 
    phi_stmt_1362_phi_mux_ack_2979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1362_ack_0, ack => outputPort_2_Daemon_CP_2845_elements(66)); -- 
    -- CP-element group 67:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1364_sample_start__ps
      -- CP-element group 67: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1364_sample_completed__ps
      -- CP-element group 67: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1364_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1364_sample_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1364_update_start__ps
      -- CP-element group 68: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1364_update_start_
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	70 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1364_update_completed__ps
      -- 
    outputPort_2_Daemon_CP_2845_elements(69) <= outputPort_2_Daemon_CP_2845_elements(70);
    -- CP-element group 70:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	69 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1364_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(70) is a control-delay.
    cp_element_70_delay: control_delay_element  generic map(name => " 70_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_2845_elements(68), ack => outputPort_2_Daemon_CP_2845_elements(70), clk => clk, reset =>reset);
    -- CP-element group 71:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_2_2_1366_sample_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(71) is bound as output of CP function.
    -- CP-element group 72:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_2_2_1366_update_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(72) is bound as output of CP function.
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: marked-predecessors 
    -- CP-element group 73: 	76 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_2_2_1366_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_2_2_1366_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_2_2_1366_Sample/rr
      -- 
    rr_3000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(73), ack => RPIPE_noblock_obuf_2_2_1366_inst_req_0); -- 
    outputPort_2_Daemon_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(71) & outputPort_2_Daemon_CP_2845_elements(76);
      gj_outputPort_2_Daemon_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: 	75 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_2_2_1366_update_start_
      -- CP-element group 74: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_2_2_1366_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_2_2_1366_Update/cr
      -- 
    cr_3005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(74), ack => RPIPE_noblock_obuf_2_2_1366_inst_req_1); -- 
    outputPort_2_Daemon_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(72) & outputPort_2_Daemon_CP_2845_elements(75);
      gj_outputPort_2_Daemon_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	74 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_2_2_1366_sample_completed__ps
      -- CP-element group 75: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_2_2_1366_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_2_2_1366_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_2_2_1366_Sample/ra
      -- 
    ra_3001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_2_1366_inst_ack_0, ack => outputPort_2_Daemon_CP_2845_elements(75)); -- 
    -- CP-element group 76:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: marked-successors 
    -- CP-element group 76: 	73 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_2_2_1366_update_completed__ps
      -- CP-element group 76: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_2_2_1366_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_2_2_1366_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_2_2_1366_Update/ca
      -- 
    ca_3006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_2_1366_inst_ack_1, ack => outputPort_2_Daemon_CP_2845_elements(76)); -- 
    -- CP-element group 77:  join  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	9 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	12 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	11 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1367_sample_start_
      -- 
    outputPort_2_Daemon_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(9) & outputPort_2_Daemon_CP_2845_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  join  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	9 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	176 
    -- CP-element group 78: 	179 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	14 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1367_update_start_
      -- 
    outputPort_2_Daemon_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(9) & outputPort_2_Daemon_CP_2845_elements(176) & outputPort_2_Daemon_CP_2845_elements(179);
      gj_outputPort_2_Daemon_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	11 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1367_sample_start__ps
      -- 
    outputPort_2_Daemon_CP_2845_elements(79) <= outputPort_2_Daemon_CP_2845_elements(11);
    -- CP-element group 80:  join  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	12 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1367_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(80) is bound as output of CP function.
    -- CP-element group 81:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	14 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1367_update_start__ps
      -- 
    outputPort_2_Daemon_CP_2845_elements(81) <= outputPort_2_Daemon_CP_2845_elements(14);
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	174 
    -- CP-element group 82: 	178 
    -- CP-element group 82: 	15 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1367_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1367_update_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(82) is bound as output of CP function.
    -- CP-element group 83:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	7 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1367_loopback_trigger
      -- 
    outputPort_2_Daemon_CP_2845_elements(83) <= outputPort_2_Daemon_CP_2845_elements(7);
    -- CP-element group 84:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1367_loopback_sample_req
      -- CP-element group 84: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1367_loopback_sample_req_ps
      -- 
    phi_stmt_1367_loopback_sample_req_3017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1367_loopback_sample_req_3017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(84), ack => phi_stmt_1367_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(84) is bound as output of CP function.
    -- CP-element group 85:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	8 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1367_entry_trigger
      -- 
    outputPort_2_Daemon_CP_2845_elements(85) <= outputPort_2_Daemon_CP_2845_elements(8);
    -- CP-element group 86:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1367_entry_sample_req
      -- CP-element group 86: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1367_entry_sample_req_ps
      -- 
    phi_stmt_1367_entry_sample_req_3020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1367_entry_sample_req_3020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(86), ack => phi_stmt_1367_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(86) is bound as output of CP function.
    -- CP-element group 87:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1367_phi_mux_ack
      -- CP-element group 87: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1367_phi_mux_ack_ps
      -- 
    phi_stmt_1367_phi_mux_ack_3023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1367_ack_0, ack => outputPort_2_Daemon_CP_2845_elements(87)); -- 
    -- CP-element group 88:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (4) 
      -- CP-element group 88: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1369_sample_start__ps
      -- CP-element group 88: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1369_sample_completed__ps
      -- CP-element group 88: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1369_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1369_sample_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1369_update_start__ps
      -- CP-element group 89: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1369_update_start_
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(89) is bound as output of CP function.
    -- CP-element group 90:  join  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	91 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1369_update_completed__ps
      -- 
    outputPort_2_Daemon_CP_2845_elements(90) <= outputPort_2_Daemon_CP_2845_elements(91);
    -- CP-element group 91:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	90 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1369_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(91) is a control-delay.
    cp_element_91_delay: control_delay_element  generic map(name => " 91_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_2845_elements(89), ack => outputPort_2_Daemon_CP_2845_elements(91), clk => clk, reset =>reset);
    -- CP-element group 92:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_3_2_1371_sample_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(92) is bound as output of CP function.
    -- CP-element group 93:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_3_2_1371_update_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(93) is bound as output of CP function.
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	97 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_3_2_1371_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_3_2_1371_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_3_2_1371_Sample/rr
      -- 
    rr_3044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(94), ack => RPIPE_noblock_obuf_3_2_1371_inst_req_0); -- 
    outputPort_2_Daemon_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(92) & outputPort_2_Daemon_CP_2845_elements(97);
      gj_outputPort_2_Daemon_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: 	96 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_3_2_1371_update_start_
      -- CP-element group 95: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_3_2_1371_Update/$entry
      -- CP-element group 95: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_3_2_1371_Update/cr
      -- 
    cr_3049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(95), ack => RPIPE_noblock_obuf_3_2_1371_inst_req_1); -- 
    outputPort_2_Daemon_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(93) & outputPort_2_Daemon_CP_2845_elements(96);
      gj_outputPort_2_Daemon_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	95 
    -- CP-element group 96:  members (4) 
      -- CP-element group 96: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_3_2_1371_sample_completed__ps
      -- CP-element group 96: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_3_2_1371_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_3_2_1371_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_3_2_1371_Sample/ra
      -- 
    ra_3045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_2_1371_inst_ack_0, ack => outputPort_2_Daemon_CP_2845_elements(96)); -- 
    -- CP-element group 97:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: marked-successors 
    -- CP-element group 97: 	94 
    -- CP-element group 97:  members (4) 
      -- CP-element group 97: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_3_2_1371_update_completed__ps
      -- CP-element group 97: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_3_2_1371_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_3_2_1371_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_3_2_1371_Update/ca
      -- 
    ca_3050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_2_1371_inst_ack_1, ack => outputPort_2_Daemon_CP_2845_elements(97)); -- 
    -- CP-element group 98:  join  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	9 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	12 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	11 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1372_sample_start_
      -- 
    outputPort_2_Daemon_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(9) & outputPort_2_Daemon_CP_2845_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  join  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	9 
    -- CP-element group 99: marked-predecessors 
    -- CP-element group 99: 	176 
    -- CP-element group 99: 	179 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	14 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1372_update_start_
      -- 
    outputPort_2_Daemon_cp_element_group_99: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_99"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(9) & outputPort_2_Daemon_CP_2845_elements(176) & outputPort_2_Daemon_CP_2845_elements(179);
      gj_outputPort_2_Daemon_cp_element_group_99 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(99), clk => clk, reset => reset); --
    end block;
    -- CP-element group 100:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	11 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1372_sample_start__ps
      -- 
    outputPort_2_Daemon_CP_2845_elements(100) <= outputPort_2_Daemon_CP_2845_elements(11);
    -- CP-element group 101:  join  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	12 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1372_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(101) is bound as output of CP function.
    -- CP-element group 102:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	14 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1372_update_start__ps
      -- 
    outputPort_2_Daemon_CP_2845_elements(102) <= outputPort_2_Daemon_CP_2845_elements(14);
    -- CP-element group 103:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	174 
    -- CP-element group 103: 	178 
    -- CP-element group 103: 	15 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1372_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1372_update_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(103) is bound as output of CP function.
    -- CP-element group 104:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	7 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1372_loopback_trigger
      -- 
    outputPort_2_Daemon_CP_2845_elements(104) <= outputPort_2_Daemon_CP_2845_elements(7);
    -- CP-element group 105:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1372_loopback_sample_req
      -- CP-element group 105: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1372_loopback_sample_req_ps
      -- 
    phi_stmt_1372_loopback_sample_req_3061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1372_loopback_sample_req_3061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(105), ack => phi_stmt_1372_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(105) is bound as output of CP function.
    -- CP-element group 106:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	8 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1372_entry_trigger
      -- 
    outputPort_2_Daemon_CP_2845_elements(106) <= outputPort_2_Daemon_CP_2845_elements(8);
    -- CP-element group 107:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1372_entry_sample_req
      -- CP-element group 107: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1372_entry_sample_req_ps
      -- 
    phi_stmt_1372_entry_sample_req_3064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1372_entry_sample_req_3064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(107), ack => phi_stmt_1372_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(107) is bound as output of CP function.
    -- CP-element group 108:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1372_phi_mux_ack
      -- CP-element group 108: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1372_phi_mux_ack_ps
      -- 
    phi_stmt_1372_phi_mux_ack_3067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1372_ack_0, ack => outputPort_2_Daemon_CP_2845_elements(108)); -- 
    -- CP-element group 109:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (4) 
      -- CP-element group 109: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1374_sample_start__ps
      -- CP-element group 109: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1374_sample_completed__ps
      -- CP-element group 109: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1374_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1374_sample_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(109) is bound as output of CP function.
    -- CP-element group 110:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1374_update_start__ps
      -- CP-element group 110: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1374_update_start_
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(110) is bound as output of CP function.
    -- CP-element group 111:  join  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1374_update_completed__ps
      -- 
    outputPort_2_Daemon_CP_2845_elements(111) <= outputPort_2_Daemon_CP_2845_elements(112);
    -- CP-element group 112:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	111 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_33_1374_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(112) is a control-delay.
    cp_element_112_delay: control_delay_element  generic map(name => " 112_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_2845_elements(110), ack => outputPort_2_Daemon_CP_2845_elements(112), clk => clk, reset =>reset);
    -- CP-element group 113:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_4_2_1376_sample_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(113) is bound as output of CP function.
    -- CP-element group 114:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_4_2_1376_update_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(114) is bound as output of CP function.
    -- CP-element group 115:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: marked-predecessors 
    -- CP-element group 115: 	118 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_4_2_1376_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_4_2_1376_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_4_2_1376_Sample/rr
      -- 
    rr_3088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(115), ack => RPIPE_noblock_obuf_4_2_1376_inst_req_0); -- 
    outputPort_2_Daemon_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(113) & outputPort_2_Daemon_CP_2845_elements(118);
      gj_outputPort_2_Daemon_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: 	117 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_4_2_1376_update_start_
      -- CP-element group 116: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_4_2_1376_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_4_2_1376_Update/cr
      -- 
    cr_3093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(116), ack => RPIPE_noblock_obuf_4_2_1376_inst_req_1); -- 
    outputPort_2_Daemon_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(114) & outputPort_2_Daemon_CP_2845_elements(117);
      gj_outputPort_2_Daemon_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	116 
    -- CP-element group 117:  members (4) 
      -- CP-element group 117: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_4_2_1376_sample_completed__ps
      -- CP-element group 117: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_4_2_1376_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_4_2_1376_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_4_2_1376_Sample/ra
      -- 
    ra_3089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_2_1376_inst_ack_0, ack => outputPort_2_Daemon_CP_2845_elements(117)); -- 
    -- CP-element group 118:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: marked-successors 
    -- CP-element group 118: 	115 
    -- CP-element group 118:  members (4) 
      -- CP-element group 118: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_4_2_1376_update_completed__ps
      -- CP-element group 118: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_4_2_1376_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_4_2_1376_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/RPIPE_noblock_obuf_4_2_1376_Update/ca
      -- 
    ca_3094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_2_1376_inst_ack_1, ack => outputPort_2_Daemon_CP_2845_elements(118)); -- 
    -- CP-element group 119:  join  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	9 
    -- CP-element group 119: marked-predecessors 
    -- CP-element group 119: 	12 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	11 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1377_sample_start_
      -- 
    outputPort_2_Daemon_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(9) & outputPort_2_Daemon_CP_2845_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  join  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	9 
    -- CP-element group 120: marked-predecessors 
    -- CP-element group 120: 	176 
    -- CP-element group 120: 	179 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	14 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1377_update_start_
      -- 
    outputPort_2_Daemon_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(9) & outputPort_2_Daemon_CP_2845_elements(176) & outputPort_2_Daemon_CP_2845_elements(179);
      gj_outputPort_2_Daemon_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	11 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1377_sample_start__ps
      -- 
    outputPort_2_Daemon_CP_2845_elements(121) <= outputPort_2_Daemon_CP_2845_elements(11);
    -- CP-element group 122:  join  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	12 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1377_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(122) is bound as output of CP function.
    -- CP-element group 123:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	14 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1377_update_start__ps
      -- 
    outputPort_2_Daemon_CP_2845_elements(123) <= outputPort_2_Daemon_CP_2845_elements(14);
    -- CP-element group 124:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	174 
    -- CP-element group 124: 	178 
    -- CP-element group 124: 	15 
    -- CP-element group 124:  members (2) 
      -- CP-element group 124: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1377_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1377_update_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(124) is bound as output of CP function.
    -- CP-element group 125:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	7 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1377_loopback_trigger
      -- 
    outputPort_2_Daemon_CP_2845_elements(125) <= outputPort_2_Daemon_CP_2845_elements(7);
    -- CP-element group 126:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1377_loopback_sample_req
      -- CP-element group 126: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1377_loopback_sample_req_ps
      -- 
    phi_stmt_1377_loopback_sample_req_3105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1377_loopback_sample_req_3105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(126), ack => phi_stmt_1377_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(126) is bound as output of CP function.
    -- CP-element group 127:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	8 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1377_entry_trigger
      -- 
    outputPort_2_Daemon_CP_2845_elements(127) <= outputPort_2_Daemon_CP_2845_elements(8);
    -- CP-element group 128:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1377_entry_sample_req
      -- CP-element group 128: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1377_entry_sample_req_ps
      -- 
    phi_stmt_1377_entry_sample_req_3108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1377_entry_sample_req_3108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(128), ack => phi_stmt_1377_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(128) is bound as output of CP function.
    -- CP-element group 129:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (2) 
      -- CP-element group 129: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1377_phi_mux_ack
      -- CP-element group 129: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1377_phi_mux_ack_ps
      -- 
    phi_stmt_1377_phi_mux_ack_3111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1377_ack_0, ack => outputPort_2_Daemon_CP_2845_elements(129)); -- 
    -- CP-element group 130:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: successors 
    -- CP-element group 130:  members (4) 
      -- CP-element group 130: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_3_1379_sample_start__ps
      -- CP-element group 130: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_3_1379_sample_completed__ps
      -- CP-element group 130: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_3_1379_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_3_1379_sample_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(130) is bound as output of CP function.
    -- CP-element group 131:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (2) 
      -- CP-element group 131: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_3_1379_update_start__ps
      -- CP-element group 131: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_3_1379_update_start_
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(131) is bound as output of CP function.
    -- CP-element group 132:  join  transition  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	133 
    -- CP-element group 132: successors 
    -- CP-element group 132:  members (1) 
      -- CP-element group 132: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_3_1379_update_completed__ps
      -- 
    outputPort_2_Daemon_CP_2845_elements(132) <= outputPort_2_Daemon_CP_2845_elements(133);
    -- CP-element group 133:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	132 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_3_1379_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(133) is a control-delay.
    cp_element_133_delay: control_delay_element  generic map(name => " 133_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_2845_elements(131), ack => outputPort_2_Daemon_CP_2845_elements(133), clk => clk, reset =>reset);
    -- CP-element group 134:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (4) 
      -- CP-element group 134: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_1380_sample_start__ps
      -- CP-element group 134: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_1380_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_1380_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_1380_Sample/req
      -- 
    req_3132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(134), ack => next_active_packet_1487_1380_buf_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(134) is bound as output of CP function.
    -- CP-element group 135:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	137 
    -- CP-element group 135:  members (4) 
      -- CP-element group 135: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_1380_update_start__ps
      -- CP-element group 135: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_1380_update_start_
      -- CP-element group 135: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_1380_Update/$entry
      -- CP-element group 135: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_1380_Update/req
      -- 
    req_3137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(135), ack => next_active_packet_1487_1380_buf_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(135) is bound as output of CP function.
    -- CP-element group 136:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (4) 
      -- CP-element group 136: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_1380_sample_completed__ps
      -- CP-element group 136: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_1380_sample_completed_
      -- CP-element group 136: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_1380_Sample/$exit
      -- CP-element group 136: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_1380_Sample/ack
      -- 
    ack_3133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_1487_1380_buf_ack_0, ack => outputPort_2_Daemon_CP_2845_elements(136)); -- 
    -- CP-element group 137:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	135 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (4) 
      -- CP-element group 137: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_1380_update_completed__ps
      -- CP-element group 137: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_1380_update_completed_
      -- CP-element group 137: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_1380_Update/$exit
      -- CP-element group 137: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_1380_Update/ack
      -- 
    ack_3138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_1487_1380_buf_ack_1, ack => outputPort_2_Daemon_CP_2845_elements(137)); -- 
    -- CP-element group 138:  join  transition  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	9 
    -- CP-element group 138: marked-predecessors 
    -- CP-element group 138: 	12 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	11 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1381_sample_start_
      -- 
    outputPort_2_Daemon_cp_element_group_138: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_138"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(9) & outputPort_2_Daemon_CP_2845_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_138 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(138), clk => clk, reset => reset); --
    end block;
    -- CP-element group 139:  join  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	9 
    -- CP-element group 139: marked-predecessors 
    -- CP-element group 139: 	142 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	14 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1381_update_start_
      -- 
    outputPort_2_Daemon_cp_element_group_139: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_139"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(9) & outputPort_2_Daemon_CP_2845_elements(142);
      gj_outputPort_2_Daemon_cp_element_group_139 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(139), clk => clk, reset => reset); --
    end block;
    -- CP-element group 140:  join  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	12 
    -- CP-element group 140:  members (1) 
      -- CP-element group 140: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1381_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(140) is bound as output of CP function.
    -- CP-element group 141:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	14 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (1) 
      -- CP-element group 141: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1381_update_start__ps
      -- 
    outputPort_2_Daemon_CP_2845_elements(141) <= outputPort_2_Daemon_CP_2845_elements(14);
    -- CP-element group 142:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	15 
    -- CP-element group 142: marked-successors 
    -- CP-element group 142: 	139 
    -- CP-element group 142:  members (2) 
      -- CP-element group 142: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1381_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1381_update_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(142) is bound as output of CP function.
    -- CP-element group 143:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	7 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1381_loopback_trigger
      -- 
    outputPort_2_Daemon_CP_2845_elements(143) <= outputPort_2_Daemon_CP_2845_elements(7);
    -- CP-element group 144:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (2) 
      -- CP-element group 144: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1381_loopback_sample_req
      -- CP-element group 144: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1381_loopback_sample_req_ps
      -- 
    phi_stmt_1381_loopback_sample_req_3149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1381_loopback_sample_req_3149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(144), ack => phi_stmt_1381_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(144) is bound as output of CP function.
    -- CP-element group 145:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	8 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (1) 
      -- CP-element group 145: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1381_entry_trigger
      -- 
    outputPort_2_Daemon_CP_2845_elements(145) <= outputPort_2_Daemon_CP_2845_elements(8);
    -- CP-element group 146:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (2) 
      -- CP-element group 146: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1381_entry_sample_req
      -- CP-element group 146: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1381_entry_sample_req_ps
      -- 
    phi_stmt_1381_entry_sample_req_3152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1381_entry_sample_req_3152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(146), ack => phi_stmt_1381_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(146) is bound as output of CP function.
    -- CP-element group 147:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (2) 
      -- CP-element group 147: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1381_phi_mux_ack
      -- CP-element group 147: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1381_phi_mux_ack_ps
      -- 
    phi_stmt_1381_phi_mux_ack_3155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1381_ack_0, ack => outputPort_2_Daemon_CP_2845_elements(147)); -- 
    -- CP-element group 148:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (4) 
      -- CP-element group 148: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_8_1383_sample_start__ps
      -- CP-element group 148: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_8_1383_sample_completed__ps
      -- CP-element group 148: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_8_1383_sample_start_
      -- CP-element group 148: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_8_1383_sample_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(148) is bound as output of CP function.
    -- CP-element group 149:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	151 
    -- CP-element group 149:  members (2) 
      -- CP-element group 149: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_8_1383_update_start__ps
      -- CP-element group 149: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_8_1383_update_start_
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(149) is bound as output of CP function.
    -- CP-element group 150:  join  transition  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	151 
    -- CP-element group 150: successors 
    -- CP-element group 150:  members (1) 
      -- CP-element group 150: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_8_1383_update_completed__ps
      -- 
    outputPort_2_Daemon_CP_2845_elements(150) <= outputPort_2_Daemon_CP_2845_elements(151);
    -- CP-element group 151:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	149 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	150 
    -- CP-element group 151:  members (1) 
      -- CP-element group 151: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_8_1383_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(151) is a control-delay.
    cp_element_151_delay: control_delay_element  generic map(name => " 151_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_2845_elements(149), ack => outputPort_2_Daemon_CP_2845_elements(151), clk => clk, reset =>reset);
    -- CP-element group 152:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (4) 
      -- CP-element group 152: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_length_1384_sample_start__ps
      -- CP-element group 152: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_length_1384_sample_start_
      -- CP-element group 152: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_length_1384_Sample/$entry
      -- CP-element group 152: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_length_1384_Sample/req
      -- 
    req_3176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(152), ack => next_active_packet_length_1532_1384_buf_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(152) is bound as output of CP function.
    -- CP-element group 153:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	155 
    -- CP-element group 153:  members (4) 
      -- CP-element group 153: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_length_1384_update_start__ps
      -- CP-element group 153: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_length_1384_update_start_
      -- CP-element group 153: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_length_1384_Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_length_1384_Update/req
      -- 
    req_3181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(153), ack => next_active_packet_length_1532_1384_buf_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(153) is bound as output of CP function.
    -- CP-element group 154:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	152 
    -- CP-element group 154: successors 
    -- CP-element group 154:  members (4) 
      -- CP-element group 154: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_length_1384_sample_completed__ps
      -- CP-element group 154: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_length_1384_sample_completed_
      -- CP-element group 154: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_length_1384_Sample/$exit
      -- CP-element group 154: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_length_1384_Sample/ack
      -- 
    ack_3177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_length_1532_1384_buf_ack_0, ack => outputPort_2_Daemon_CP_2845_elements(154)); -- 
    -- CP-element group 155:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	153 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (4) 
      -- CP-element group 155: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_length_1384_update_completed__ps
      -- CP-element group 155: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_length_1384_update_completed_
      -- CP-element group 155: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_length_1384_Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_active_packet_length_1384_Update/ack
      -- 
    ack_3182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_length_1532_1384_buf_ack_1, ack => outputPort_2_Daemon_CP_2845_elements(155)); -- 
    -- CP-element group 156:  join  transition  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	9 
    -- CP-element group 156: marked-predecessors 
    -- CP-element group 156: 	12 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	11 
    -- CP-element group 156:  members (1) 
      -- CP-element group 156: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1385_sample_start_
      -- 
    outputPort_2_Daemon_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(9) & outputPort_2_Daemon_CP_2845_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  join  transition  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	9 
    -- CP-element group 157: marked-predecessors 
    -- CP-element group 157: 	176 
    -- CP-element group 157: 	179 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	14 
    -- CP-element group 157:  members (1) 
      -- CP-element group 157: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1385_update_start_
      -- 
    outputPort_2_Daemon_cp_element_group_157: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_157"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(9) & outputPort_2_Daemon_CP_2845_elements(176) & outputPort_2_Daemon_CP_2845_elements(179);
      gj_outputPort_2_Daemon_cp_element_group_157 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(157), clk => clk, reset => reset); --
    end block;
    -- CP-element group 158:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	11 
    -- CP-element group 158: successors 
    -- CP-element group 158:  members (1) 
      -- CP-element group 158: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1385_sample_start__ps
      -- 
    outputPort_2_Daemon_CP_2845_elements(158) <= outputPort_2_Daemon_CP_2845_elements(11);
    -- CP-element group 159:  join  transition  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	12 
    -- CP-element group 159:  members (1) 
      -- CP-element group 159: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1385_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(159) is bound as output of CP function.
    -- CP-element group 160:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	174 
    -- CP-element group 160: 	178 
    -- CP-element group 160: 	15 
    -- CP-element group 160:  members (2) 
      -- CP-element group 160: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1385_update_completed_
      -- CP-element group 160: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1385_update_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(160) is bound as output of CP function.
    -- CP-element group 161:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	7 
    -- CP-element group 161: successors 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1385_loopback_trigger
      -- 
    outputPort_2_Daemon_CP_2845_elements(161) <= outputPort_2_Daemon_CP_2845_elements(7);
    -- CP-element group 162:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (2) 
      -- CP-element group 162: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1385_loopback_sample_req_ps
      -- CP-element group 162: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1385_loopback_sample_req
      -- 
    phi_stmt_1385_loopback_sample_req_3193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1385_loopback_sample_req_3193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(162), ack => phi_stmt_1385_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(162) is bound as output of CP function.
    -- CP-element group 163:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	8 
    -- CP-element group 163: successors 
    -- CP-element group 163:  members (1) 
      -- CP-element group 163: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1385_entry_trigger
      -- 
    outputPort_2_Daemon_CP_2845_elements(163) <= outputPort_2_Daemon_CP_2845_elements(8);
    -- CP-element group 164:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (2) 
      -- CP-element group 164: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1385_entry_sample_req_ps
      -- CP-element group 164: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1385_entry_sample_req
      -- 
    phi_stmt_1385_entry_sample_req_3196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1385_entry_sample_req_3196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(164), ack => phi_stmt_1385_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(164) is bound as output of CP function.
    -- CP-element group 165:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: successors 
    -- CP-element group 165:  members (2) 
      -- CP-element group 165: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1385_phi_mux_ack_ps
      -- CP-element group 165: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/phi_stmt_1385_phi_mux_ack
      -- 
    phi_stmt_1385_phi_mux_ack_3199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1385_ack_0, ack => outputPort_2_Daemon_CP_2845_elements(165)); -- 
    -- CP-element group 166:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: successors 
    -- CP-element group 166:  members (4) 
      -- CP-element group 166: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_2_1387_sample_start__ps
      -- CP-element group 166: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_2_1387_sample_start_
      -- CP-element group 166: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_2_1387_sample_completed_
      -- CP-element group 166: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_2_1387_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(166) is bound as output of CP function.
    -- CP-element group 167:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (2) 
      -- CP-element group 167: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_2_1387_update_start__ps
      -- CP-element group 167: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_2_1387_update_start_
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(167) is bound as output of CP function.
    -- CP-element group 168:  join  transition  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	169 
    -- CP-element group 168: successors 
    -- CP-element group 168:  members (1) 
      -- CP-element group 168: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_2_1387_update_completed__ps
      -- 
    outputPort_2_Daemon_CP_2845_elements(168) <= outputPort_2_Daemon_CP_2845_elements(169);
    -- CP-element group 169:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	168 
    -- CP-element group 169:  members (1) 
      -- CP-element group 169: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_ZERO_2_1387_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(169) is a control-delay.
    cp_element_169_delay: control_delay_element  generic map(name => " 169_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_2845_elements(167), ack => outputPort_2_Daemon_CP_2845_elements(169), clk => clk, reset =>reset);
    -- CP-element group 170:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	172 
    -- CP-element group 170:  members (4) 
      -- CP-element group 170: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_priority_index_1388_sample_start__ps
      -- CP-element group 170: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_priority_index_1388_sample_start_
      -- CP-element group 170: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_priority_index_1388_Sample/req
      -- CP-element group 170: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_priority_index_1388_Sample/$entry
      -- 
    req_3220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(170), ack => next_priority_index_1487_1388_buf_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(170) is bound as output of CP function.
    -- CP-element group 171:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (4) 
      -- CP-element group 171: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_priority_index_1388_update_start__ps
      -- CP-element group 171: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_priority_index_1388_Update/req
      -- CP-element group 171: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_priority_index_1388_Update/$entry
      -- CP-element group 171: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_priority_index_1388_update_start_
      -- 
    req_3225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(171), ack => next_priority_index_1487_1388_buf_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(171) is bound as output of CP function.
    -- CP-element group 172:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	170 
    -- CP-element group 172: successors 
    -- CP-element group 172:  members (4) 
      -- CP-element group 172: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_priority_index_1388_sample_completed__ps
      -- CP-element group 172: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_priority_index_1388_Sample/ack
      -- CP-element group 172: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_priority_index_1388_Sample/$exit
      -- CP-element group 172: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_priority_index_1388_sample_completed_
      -- 
    ack_3221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_priority_index_1487_1388_buf_ack_0, ack => outputPort_2_Daemon_CP_2845_elements(172)); -- 
    -- CP-element group 173:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: successors 
    -- CP-element group 173:  members (4) 
      -- CP-element group 173: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_priority_index_1388_update_completed__ps
      -- CP-element group 173: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_priority_index_1388_Update/ack
      -- CP-element group 173: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_priority_index_1388_Update/$exit
      -- CP-element group 173: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/R_next_priority_index_1388_update_completed_
      -- 
    ack_3226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_priority_index_1487_1388_buf_ack_1, ack => outputPort_2_Daemon_CP_2845_elements(173)); -- 
    -- CP-element group 174:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	160 
    -- CP-element group 174: 	21 
    -- CP-element group 174: 	40 
    -- CP-element group 174: 	61 
    -- CP-element group 174: 	82 
    -- CP-element group 174: 	103 
    -- CP-element group 174: 	124 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	176 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/call_stmt_1416_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/call_stmt_1416_Sample/crr
      -- CP-element group 174: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/call_stmt_1416_Sample/$entry
      -- 
    crr_3235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(174), ack => call_stmt_1416_call_req_0); -- 
    outputPort_2_Daemon_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(160) & outputPort_2_Daemon_CP_2845_elements(21) & outputPort_2_Daemon_CP_2845_elements(40) & outputPort_2_Daemon_CP_2845_elements(61) & outputPort_2_Daemon_CP_2845_elements(82) & outputPort_2_Daemon_CP_2845_elements(103) & outputPort_2_Daemon_CP_2845_elements(124);
      gj_outputPort_2_Daemon_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: marked-predecessors 
    -- CP-element group 175: 	177 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	177 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/call_stmt_1416_Update/ccr
      -- CP-element group 175: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/call_stmt_1416_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/call_stmt_1416_update_start_
      -- 
    ccr_3240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(175), ack => call_stmt_1416_call_req_1); -- 
    outputPort_2_Daemon_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= outputPort_2_Daemon_CP_2845_elements(177);
      gj_outputPort_2_Daemon_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	174 
    -- CP-element group 176: successors 
    -- CP-element group 176: marked-successors 
    -- CP-element group 176: 	157 
    -- CP-element group 176: 	17 
    -- CP-element group 176: 	36 
    -- CP-element group 176: 	57 
    -- CP-element group 176: 	78 
    -- CP-element group 176: 	99 
    -- CP-element group 176: 	120 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/call_stmt_1416_Sample/cra
      -- CP-element group 176: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/call_stmt_1416_Sample/$exit
      -- CP-element group 176: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/call_stmt_1416_sample_completed_
      -- 
    cra_3236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1416_call_ack_0, ack => outputPort_2_Daemon_CP_2845_elements(176)); -- 
    -- CP-element group 177:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	182 
    -- CP-element group 177: marked-successors 
    -- CP-element group 177: 	175 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/call_stmt_1416_Update/$exit
      -- CP-element group 177: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/call_stmt_1416_Update/cca
      -- CP-element group 177: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/call_stmt_1416_update_completed_
      -- 
    cca_3241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1416_call_ack_1, ack => outputPort_2_Daemon_CP_2845_elements(177)); -- 
    -- CP-element group 178:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	160 
    -- CP-element group 178: 	21 
    -- CP-element group 178: 	40 
    -- CP-element group 178: 	61 
    -- CP-element group 178: 	82 
    -- CP-element group 178: 	103 
    -- CP-element group 178: 	124 
    -- CP-element group 178: marked-predecessors 
    -- CP-element group 178: 	180 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/WPIPE_out_data_2_1641_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/WPIPE_out_data_2_1641_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/WPIPE_out_data_2_1641_Sample/req
      -- 
    req_3249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(178), ack => WPIPE_out_data_2_1641_inst_req_0); -- 
    outputPort_2_Daemon_cp_element_group_178: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_178"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(160) & outputPort_2_Daemon_CP_2845_elements(21) & outputPort_2_Daemon_CP_2845_elements(40) & outputPort_2_Daemon_CP_2845_elements(61) & outputPort_2_Daemon_CP_2845_elements(82) & outputPort_2_Daemon_CP_2845_elements(103) & outputPort_2_Daemon_CP_2845_elements(124) & outputPort_2_Daemon_CP_2845_elements(180);
      gj_outputPort_2_Daemon_cp_element_group_178 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(178), clk => clk, reset => reset); --
    end block;
    -- CP-element group 179:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179: marked-successors 
    -- CP-element group 179: 	157 
    -- CP-element group 179: 	17 
    -- CP-element group 179: 	36 
    -- CP-element group 179: 	57 
    -- CP-element group 179: 	78 
    -- CP-element group 179: 	99 
    -- CP-element group 179: 	120 
    -- CP-element group 179:  members (6) 
      -- CP-element group 179: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/WPIPE_out_data_2_1641_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/WPIPE_out_data_2_1641_update_start_
      -- CP-element group 179: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/WPIPE_out_data_2_1641_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/WPIPE_out_data_2_1641_Sample/ack
      -- CP-element group 179: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/WPIPE_out_data_2_1641_Update/$entry
      -- CP-element group 179: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/WPIPE_out_data_2_1641_Update/req
      -- 
    ack_3250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_2_1641_inst_ack_0, ack => outputPort_2_Daemon_CP_2845_elements(179)); -- 
    req_3254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_2845_elements(179), ack => WPIPE_out_data_2_1641_inst_req_1); -- 
    -- CP-element group 180:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	182 
    -- CP-element group 180: marked-successors 
    -- CP-element group 180: 	178 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/WPIPE_out_data_2_1641_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/WPIPE_out_data_2_1641_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/WPIPE_out_data_2_1641_Update/ack
      -- 
    ack_3255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_2_1641_inst_ack_1, ack => outputPort_2_Daemon_CP_2845_elements(180)); -- 
    -- CP-element group 181:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	9 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	10 
    -- CP-element group 181:  members (1) 
      -- CP-element group 181: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group outputPort_2_Daemon_CP_2845_elements(181) is a control-delay.
    cp_element_181_delay: control_delay_element  generic map(name => " 181_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_2845_elements(9), ack => outputPort_2_Daemon_CP_2845_elements(181), clk => clk, reset =>reset);
    -- CP-element group 182:  join  transition  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	180 
    -- CP-element group 182: 	177 
    -- CP-element group 182: 	12 
    -- CP-element group 182: 	13 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	6 
    -- CP-element group 182:  members (1) 
      -- CP-element group 182: 	 branch_block_stmt_1350/do_while_stmt_1351/do_while_stmt_1351_loop_body/$exit
      -- 
    outputPort_2_Daemon_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 7,2 => 7,3 => 7);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_2845_elements(180) & outputPort_2_Daemon_CP_2845_elements(177) & outputPort_2_Daemon_CP_2845_elements(12) & outputPort_2_Daemon_CP_2845_elements(13);
      gj_outputPort_2_Daemon_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  transition  input  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	5 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (2) 
      -- CP-element group 183: 	 branch_block_stmt_1350/do_while_stmt_1351/loop_exit/$exit
      -- CP-element group 183: 	 branch_block_stmt_1350/do_while_stmt_1351/loop_exit/ack
      -- 
    ack_3260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1351_branch_ack_0, ack => outputPort_2_Daemon_CP_2845_elements(183)); -- 
    -- CP-element group 184:  transition  input  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	5 
    -- CP-element group 184: successors 
    -- CP-element group 184:  members (2) 
      -- CP-element group 184: 	 branch_block_stmt_1350/do_while_stmt_1351/loop_taken/$exit
      -- CP-element group 184: 	 branch_block_stmt_1350/do_while_stmt_1351/loop_taken/ack
      -- 
    ack_3264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1351_branch_ack_1, ack => outputPort_2_Daemon_CP_2845_elements(184)); -- 
    -- CP-element group 185:  transition  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	3 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	1 
    -- CP-element group 185:  members (1) 
      -- CP-element group 185: 	 branch_block_stmt_1350/do_while_stmt_1351/$exit
      -- 
    outputPort_2_Daemon_CP_2845_elements(185) <= outputPort_2_Daemon_CP_2845_elements(3);
    outputPort_2_Daemon_do_while_stmt_1351_terminator_3265: loop_terminator -- 
      generic map (name => " outputPort_2_Daemon_do_while_stmt_1351_terminator_3265", max_iterations_in_flight =>7) 
      port map(loop_body_exit => outputPort_2_Daemon_CP_2845_elements(6),loop_continue => outputPort_2_Daemon_CP_2845_elements(184),loop_terminate => outputPort_2_Daemon_CP_2845_elements(183),loop_back => outputPort_2_Daemon_CP_2845_elements(4),loop_exit => outputPort_2_Daemon_CP_2845_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1353_phi_seq_2919_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_2_Daemon_CP_2845_elements(24);
      outputPort_2_Daemon_CP_2845_elements(27)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_2_Daemon_CP_2845_elements(27);
      outputPort_2_Daemon_CP_2845_elements(28)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_2_Daemon_CP_2845_elements(29);
      outputPort_2_Daemon_CP_2845_elements(25) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_2_Daemon_CP_2845_elements(22);
      outputPort_2_Daemon_CP_2845_elements(31)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_2_Daemon_CP_2845_elements(33);
      outputPort_2_Daemon_CP_2845_elements(32)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_2_Daemon_CP_2845_elements(34);
      outputPort_2_Daemon_CP_2845_elements(23) <= phi_mux_reqs(1);
      phi_stmt_1353_phi_seq_2919 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1353_phi_seq_2919") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_2_Daemon_CP_2845_elements(18), 
          phi_sample_ack => outputPort_2_Daemon_CP_2845_elements(19), 
          phi_update_req => outputPort_2_Daemon_CP_2845_elements(20), 
          phi_update_ack => outputPort_2_Daemon_CP_2845_elements(21), 
          phi_mux_ack => outputPort_2_Daemon_CP_2845_elements(26), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1357_phi_seq_2963_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_2_Daemon_CP_2845_elements(43);
      outputPort_2_Daemon_CP_2845_elements(46)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_2_Daemon_CP_2845_elements(46);
      outputPort_2_Daemon_CP_2845_elements(47)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_2_Daemon_CP_2845_elements(48);
      outputPort_2_Daemon_CP_2845_elements(44) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_2_Daemon_CP_2845_elements(41);
      outputPort_2_Daemon_CP_2845_elements(50)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_2_Daemon_CP_2845_elements(54);
      outputPort_2_Daemon_CP_2845_elements(51)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_2_Daemon_CP_2845_elements(55);
      outputPort_2_Daemon_CP_2845_elements(42) <= phi_mux_reqs(1);
      phi_stmt_1357_phi_seq_2963 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1357_phi_seq_2963") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_2_Daemon_CP_2845_elements(37), 
          phi_sample_ack => outputPort_2_Daemon_CP_2845_elements(38), 
          phi_update_req => outputPort_2_Daemon_CP_2845_elements(39), 
          phi_update_ack => outputPort_2_Daemon_CP_2845_elements(40), 
          phi_mux_ack => outputPort_2_Daemon_CP_2845_elements(45), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1362_phi_seq_3007_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_2_Daemon_CP_2845_elements(64);
      outputPort_2_Daemon_CP_2845_elements(67)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_2_Daemon_CP_2845_elements(67);
      outputPort_2_Daemon_CP_2845_elements(68)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_2_Daemon_CP_2845_elements(69);
      outputPort_2_Daemon_CP_2845_elements(65) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_2_Daemon_CP_2845_elements(62);
      outputPort_2_Daemon_CP_2845_elements(71)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_2_Daemon_CP_2845_elements(75);
      outputPort_2_Daemon_CP_2845_elements(72)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_2_Daemon_CP_2845_elements(76);
      outputPort_2_Daemon_CP_2845_elements(63) <= phi_mux_reqs(1);
      phi_stmt_1362_phi_seq_3007 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1362_phi_seq_3007") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_2_Daemon_CP_2845_elements(58), 
          phi_sample_ack => outputPort_2_Daemon_CP_2845_elements(59), 
          phi_update_req => outputPort_2_Daemon_CP_2845_elements(60), 
          phi_update_ack => outputPort_2_Daemon_CP_2845_elements(61), 
          phi_mux_ack => outputPort_2_Daemon_CP_2845_elements(66), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1367_phi_seq_3051_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_2_Daemon_CP_2845_elements(85);
      outputPort_2_Daemon_CP_2845_elements(88)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_2_Daemon_CP_2845_elements(88);
      outputPort_2_Daemon_CP_2845_elements(89)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_2_Daemon_CP_2845_elements(90);
      outputPort_2_Daemon_CP_2845_elements(86) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_2_Daemon_CP_2845_elements(83);
      outputPort_2_Daemon_CP_2845_elements(92)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_2_Daemon_CP_2845_elements(96);
      outputPort_2_Daemon_CP_2845_elements(93)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_2_Daemon_CP_2845_elements(97);
      outputPort_2_Daemon_CP_2845_elements(84) <= phi_mux_reqs(1);
      phi_stmt_1367_phi_seq_3051 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1367_phi_seq_3051") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_2_Daemon_CP_2845_elements(79), 
          phi_sample_ack => outputPort_2_Daemon_CP_2845_elements(80), 
          phi_update_req => outputPort_2_Daemon_CP_2845_elements(81), 
          phi_update_ack => outputPort_2_Daemon_CP_2845_elements(82), 
          phi_mux_ack => outputPort_2_Daemon_CP_2845_elements(87), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1372_phi_seq_3095_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_2_Daemon_CP_2845_elements(106);
      outputPort_2_Daemon_CP_2845_elements(109)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_2_Daemon_CP_2845_elements(109);
      outputPort_2_Daemon_CP_2845_elements(110)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_2_Daemon_CP_2845_elements(111);
      outputPort_2_Daemon_CP_2845_elements(107) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_2_Daemon_CP_2845_elements(104);
      outputPort_2_Daemon_CP_2845_elements(113)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_2_Daemon_CP_2845_elements(117);
      outputPort_2_Daemon_CP_2845_elements(114)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_2_Daemon_CP_2845_elements(118);
      outputPort_2_Daemon_CP_2845_elements(105) <= phi_mux_reqs(1);
      phi_stmt_1372_phi_seq_3095 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1372_phi_seq_3095") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_2_Daemon_CP_2845_elements(100), 
          phi_sample_ack => outputPort_2_Daemon_CP_2845_elements(101), 
          phi_update_req => outputPort_2_Daemon_CP_2845_elements(102), 
          phi_update_ack => outputPort_2_Daemon_CP_2845_elements(103), 
          phi_mux_ack => outputPort_2_Daemon_CP_2845_elements(108), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1377_phi_seq_3139_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_2_Daemon_CP_2845_elements(127);
      outputPort_2_Daemon_CP_2845_elements(130)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_2_Daemon_CP_2845_elements(130);
      outputPort_2_Daemon_CP_2845_elements(131)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_2_Daemon_CP_2845_elements(132);
      outputPort_2_Daemon_CP_2845_elements(128) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_2_Daemon_CP_2845_elements(125);
      outputPort_2_Daemon_CP_2845_elements(134)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_2_Daemon_CP_2845_elements(136);
      outputPort_2_Daemon_CP_2845_elements(135)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_2_Daemon_CP_2845_elements(137);
      outputPort_2_Daemon_CP_2845_elements(126) <= phi_mux_reqs(1);
      phi_stmt_1377_phi_seq_3139 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1377_phi_seq_3139") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_2_Daemon_CP_2845_elements(121), 
          phi_sample_ack => outputPort_2_Daemon_CP_2845_elements(122), 
          phi_update_req => outputPort_2_Daemon_CP_2845_elements(123), 
          phi_update_ack => outputPort_2_Daemon_CP_2845_elements(124), 
          phi_mux_ack => outputPort_2_Daemon_CP_2845_elements(129), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1381_phi_seq_3183_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_2_Daemon_CP_2845_elements(145);
      outputPort_2_Daemon_CP_2845_elements(148)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_2_Daemon_CP_2845_elements(148);
      outputPort_2_Daemon_CP_2845_elements(149)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_2_Daemon_CP_2845_elements(150);
      outputPort_2_Daemon_CP_2845_elements(146) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_2_Daemon_CP_2845_elements(143);
      outputPort_2_Daemon_CP_2845_elements(152)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_2_Daemon_CP_2845_elements(154);
      outputPort_2_Daemon_CP_2845_elements(153)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_2_Daemon_CP_2845_elements(155);
      outputPort_2_Daemon_CP_2845_elements(144) <= phi_mux_reqs(1);
      phi_stmt_1381_phi_seq_3183 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1381_phi_seq_3183") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_2_Daemon_CP_2845_elements(11), 
          phi_sample_ack => outputPort_2_Daemon_CP_2845_elements(140), 
          phi_update_req => outputPort_2_Daemon_CP_2845_elements(141), 
          phi_update_ack => outputPort_2_Daemon_CP_2845_elements(142), 
          phi_mux_ack => outputPort_2_Daemon_CP_2845_elements(147), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1385_phi_seq_3227_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_2_Daemon_CP_2845_elements(163);
      outputPort_2_Daemon_CP_2845_elements(166)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_2_Daemon_CP_2845_elements(166);
      outputPort_2_Daemon_CP_2845_elements(167)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_2_Daemon_CP_2845_elements(168);
      outputPort_2_Daemon_CP_2845_elements(164) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_2_Daemon_CP_2845_elements(161);
      outputPort_2_Daemon_CP_2845_elements(170)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_2_Daemon_CP_2845_elements(172);
      outputPort_2_Daemon_CP_2845_elements(171)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_2_Daemon_CP_2845_elements(173);
      outputPort_2_Daemon_CP_2845_elements(162) <= phi_mux_reqs(1);
      phi_stmt_1385_phi_seq_3227 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1385_phi_seq_3227") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_2_Daemon_CP_2845_elements(158), 
          phi_sample_ack => outputPort_2_Daemon_CP_2845_elements(159), 
          phi_update_req => outputPort_2_Daemon_CP_2845_elements(14), 
          phi_update_ack => outputPort_2_Daemon_CP_2845_elements(160), 
          phi_mux_ack => outputPort_2_Daemon_CP_2845_elements(165), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_2870_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= outputPort_2_Daemon_CP_2845_elements(7);
        preds(1)  <= outputPort_2_Daemon_CP_2845_elements(8);
        entry_tmerge_2870 : transition_merge -- 
          generic map(name => " entry_tmerge_2870")
          port map (preds => preds, symbol_out => outputPort_2_Daemon_CP_2845_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal EQ_u3_u1_1452_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1458_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1465_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1471_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1501_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1508_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1516_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1523_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1551_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1559_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1567_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1575_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1581_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1588_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1596_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1603_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1614_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1620_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1627_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1633_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_1494_wire : std_logic_vector(0 downto 0);
    signal MUX_1394_wire : std_logic_vector(7 downto 0);
    signal MUX_1398_wire : std_logic_vector(7 downto 0);
    signal MUX_1403_wire : std_logic_vector(7 downto 0);
    signal MUX_1407_wire : std_logic_vector(7 downto 0);
    signal MUX_1455_wire : std_logic_vector(0 downto 0);
    signal MUX_1461_wire : std_logic_vector(0 downto 0);
    signal MUX_1468_wire : std_logic_vector(0 downto 0);
    signal MUX_1474_wire : std_logic_vector(0 downto 0);
    signal MUX_1505_wire : std_logic_vector(7 downto 0);
    signal MUX_1512_wire : std_logic_vector(7 downto 0);
    signal MUX_1520_wire : std_logic_vector(7 downto 0);
    signal MUX_1527_wire : std_logic_vector(7 downto 0);
    signal MUX_1543_wire : std_logic_vector(7 downto 0);
    signal MUX_1585_wire : std_logic_vector(31 downto 0);
    signal MUX_1592_wire : std_logic_vector(31 downto 0);
    signal MUX_1600_wire : std_logic_vector(31 downto 0);
    signal MUX_1607_wire : std_logic_vector(31 downto 0);
    signal MUX_1617_wire : std_logic_vector(0 downto 0);
    signal MUX_1623_wire : std_logic_vector(0 downto 0);
    signal MUX_1630_wire : std_logic_vector(0 downto 0);
    signal MUX_1636_wire : std_logic_vector(0 downto 0);
    signal NEQ_u3_u1_1491_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1548_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1556_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1564_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1572_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1462_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1475_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1624_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1637_wire : std_logic_vector(0 downto 0);
    signal OR_u32_u32_1593_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_1608_wire : std_logic_vector(31 downto 0);
    signal OR_u8_u8_1399_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_1408_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_1513_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_1528_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_1529_wire : std_logic_vector(7 downto 0);
    signal RPIPE_noblock_obuf_1_2_1361_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_2_2_1366_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_3_2_1371_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_4_2_1376_wire : std_logic_vector(32 downto 0);
    signal R_ZERO_2_1387_wire_constant : std_logic_vector(1 downto 0);
    signal R_ZERO_33_1359_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1364_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1369_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1374_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_3_1379_wire_constant : std_logic_vector(2 downto 0);
    signal R_ZERO_8_1355_wire_constant : std_logic_vector(7 downto 0);
    signal R_ZERO_8_1383_wire_constant : std_logic_vector(7 downto 0);
    signal SUB_u8_u8_1537_wire : std_logic_vector(7 downto 0);
    signal SUB_u8_u8_1541_wire : std_logic_vector(7 downto 0);
    signal active_packet_1377 : std_logic_vector(2 downto 0);
    signal active_packet_length_1381 : std_logic_vector(7 downto 0);
    signal continue_1416 : std_logic_vector(0 downto 0);
    signal data_to_out_1610 : std_logic_vector(31 downto 0);
    signal down_counter_1353 : std_logic_vector(7 downto 0);
    signal konst_1392_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1393_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1396_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1397_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1401_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1402_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1405_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1406_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1412_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1419_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1424_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1429_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1434_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1451_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1454_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1457_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1460_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1464_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1467_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1470_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1473_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1490_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1493_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1500_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1504_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1507_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1511_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1515_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1519_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1522_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1526_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1536_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1540_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1550_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1558_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1566_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1574_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1580_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1584_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1587_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1591_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1595_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1599_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1602_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1606_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1613_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1616_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1619_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1622_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1626_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1629_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1632_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1635_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1654_wire_constant : std_logic_vector(0 downto 0);
    signal next_active_packet_1487 : std_logic_vector(2 downto 0);
    signal next_active_packet_1487_1380_buffered : std_logic_vector(2 downto 0);
    signal next_active_packet_length_1532 : std_logic_vector(7 downto 0);
    signal next_active_packet_length_1532_1384_buffered : std_logic_vector(7 downto 0);
    signal next_down_counter_1545 : std_logic_vector(7 downto 0);
    signal next_down_counter_1545_1356_buffered : std_logic_vector(7 downto 0);
    signal next_priority_index_1487 : std_logic_vector(1 downto 0);
    signal next_priority_index_1487_1388_buffered : std_logic_vector(1 downto 0);
    signal p1_valid_1421 : std_logic_vector(0 downto 0);
    signal p2_valid_1426 : std_logic_vector(0 downto 0);
    signal p3_valid_1431 : std_logic_vector(0 downto 0);
    signal p4_valid_1436 : std_logic_vector(0 downto 0);
    signal pkt_1_e_word_1357 : std_logic_vector(32 downto 0);
    signal pkt_2_e_word_1362 : std_logic_vector(32 downto 0);
    signal pkt_3_e_word_1367 : std_logic_vector(32 downto 0);
    signal pkt_4_e_word_1372 : std_logic_vector(32 downto 0);
    signal priority_index_1385 : std_logic_vector(1 downto 0);
    signal read_from_1_1553 : std_logic_vector(0 downto 0);
    signal read_from_2_1561 : std_logic_vector(0 downto 0);
    signal read_from_3_1569 : std_logic_vector(0 downto 0);
    signal read_from_4_1577 : std_logic_vector(0 downto 0);
    signal send_flag_1639 : std_logic_vector(0 downto 0);
    signal senderPort_1410 : std_logic_vector(7 downto 0);
    signal slice_1503_wire : std_logic_vector(7 downto 0);
    signal slice_1510_wire : std_logic_vector(7 downto 0);
    signal slice_1518_wire : std_logic_vector(7 downto 0);
    signal slice_1525_wire : std_logic_vector(7 downto 0);
    signal slice_1583_wire : std_logic_vector(31 downto 0);
    signal slice_1590_wire : std_logic_vector(31 downto 0);
    signal slice_1598_wire : std_logic_vector(31 downto 0);
    signal slice_1605_wire : std_logic_vector(31 downto 0);
    signal started_new_packet_1496 : std_logic_vector(0 downto 0);
    signal type_cast_1414_wire_constant : std_logic_vector(0 downto 0);
    signal valid_active_pkt_word_read_1477 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_ZERO_2_1387_wire_constant <= "00";
    R_ZERO_33_1359_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1364_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1369_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1374_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_3_1379_wire_constant <= "000";
    R_ZERO_8_1355_wire_constant <= "00000000";
    R_ZERO_8_1383_wire_constant <= "00000000";
    konst_1392_wire_constant <= "00000000";
    konst_1393_wire_constant <= "00000000";
    konst_1396_wire_constant <= "00000001";
    konst_1397_wire_constant <= "00000000";
    konst_1401_wire_constant <= "00000010";
    konst_1402_wire_constant <= "00000000";
    konst_1405_wire_constant <= "00000011";
    konst_1406_wire_constant <= "00000000";
    konst_1412_wire_constant <= "00000001";
    konst_1419_wire_constant <= "000000000000000000000000000100000";
    konst_1424_wire_constant <= "000000000000000000000000000100000";
    konst_1429_wire_constant <= "000000000000000000000000000100000";
    konst_1434_wire_constant <= "000000000000000000000000000100000";
    konst_1451_wire_constant <= "001";
    konst_1454_wire_constant <= "0";
    konst_1457_wire_constant <= "010";
    konst_1460_wire_constant <= "0";
    konst_1464_wire_constant <= "011";
    konst_1467_wire_constant <= "0";
    konst_1470_wire_constant <= "100";
    konst_1473_wire_constant <= "0";
    konst_1490_wire_constant <= "000";
    konst_1493_wire_constant <= "00000000";
    konst_1500_wire_constant <= "001";
    konst_1504_wire_constant <= "00000000";
    konst_1507_wire_constant <= "010";
    konst_1511_wire_constant <= "00000000";
    konst_1515_wire_constant <= "011";
    konst_1519_wire_constant <= "00000000";
    konst_1522_wire_constant <= "100";
    konst_1526_wire_constant <= "00000000";
    konst_1536_wire_constant <= "00000001";
    konst_1540_wire_constant <= "00000001";
    konst_1550_wire_constant <= "001";
    konst_1558_wire_constant <= "010";
    konst_1566_wire_constant <= "011";
    konst_1574_wire_constant <= "100";
    konst_1580_wire_constant <= "001";
    konst_1584_wire_constant <= "00000000000000000000000000000000";
    konst_1587_wire_constant <= "010";
    konst_1591_wire_constant <= "00000000000000000000000000000000";
    konst_1595_wire_constant <= "011";
    konst_1599_wire_constant <= "00000000000000000000000000000000";
    konst_1602_wire_constant <= "100";
    konst_1606_wire_constant <= "00000000000000000000000000000000";
    konst_1613_wire_constant <= "001";
    konst_1616_wire_constant <= "0";
    konst_1619_wire_constant <= "010";
    konst_1622_wire_constant <= "0";
    konst_1626_wire_constant <= "011";
    konst_1629_wire_constant <= "0";
    konst_1632_wire_constant <= "100";
    konst_1635_wire_constant <= "0";
    konst_1654_wire_constant <= "1";
    type_cast_1414_wire_constant <= "0";
    phi_stmt_1353: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_8_1355_wire_constant & next_down_counter_1545_1356_buffered;
      req <= phi_stmt_1353_req_0 & phi_stmt_1353_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1353",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1353_ack_0,
          idata => idata,
          odata => down_counter_1353,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1353
    phi_stmt_1357: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1359_wire_constant & RPIPE_noblock_obuf_1_2_1361_wire;
      req <= phi_stmt_1357_req_0 & phi_stmt_1357_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1357",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1357_ack_0,
          idata => idata,
          odata => pkt_1_e_word_1357,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1357
    phi_stmt_1362: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1364_wire_constant & RPIPE_noblock_obuf_2_2_1366_wire;
      req <= phi_stmt_1362_req_0 & phi_stmt_1362_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1362",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1362_ack_0,
          idata => idata,
          odata => pkt_2_e_word_1362,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1362
    phi_stmt_1367: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1369_wire_constant & RPIPE_noblock_obuf_3_2_1371_wire;
      req <= phi_stmt_1367_req_0 & phi_stmt_1367_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1367",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1367_ack_0,
          idata => idata,
          odata => pkt_3_e_word_1367,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1367
    phi_stmt_1372: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1374_wire_constant & RPIPE_noblock_obuf_4_2_1376_wire;
      req <= phi_stmt_1372_req_0 & phi_stmt_1372_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1372",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1372_ack_0,
          idata => idata,
          odata => pkt_4_e_word_1372,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1372
    phi_stmt_1377: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_3_1379_wire_constant & next_active_packet_1487_1380_buffered;
      req <= phi_stmt_1377_req_0 & phi_stmt_1377_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1377",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1377_ack_0,
          idata => idata,
          odata => active_packet_1377,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1377
    phi_stmt_1381: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_8_1383_wire_constant & next_active_packet_length_1532_1384_buffered;
      req <= phi_stmt_1381_req_0 & phi_stmt_1381_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1381",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1381_ack_0,
          idata => idata,
          odata => active_packet_length_1381,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1381
    phi_stmt_1385: Block -- phi operator 
      signal idata: std_logic_vector(3 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_2_1387_wire_constant & next_priority_index_1487_1388_buffered;
      req <= phi_stmt_1385_req_0 & phi_stmt_1385_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1385",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 2) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1385_ack_0,
          idata => idata,
          odata => priority_index_1385,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1385
    -- flow-through select operator MUX_1394_inst
    MUX_1394_wire <= konst_1392_wire_constant when (read_from_1_1553(0) /=  '0') else konst_1393_wire_constant;
    -- flow-through select operator MUX_1398_inst
    MUX_1398_wire <= konst_1396_wire_constant when (read_from_2_1561(0) /=  '0') else konst_1397_wire_constant;
    -- flow-through select operator MUX_1403_inst
    MUX_1403_wire <= konst_1401_wire_constant when (read_from_3_1569(0) /=  '0') else konst_1402_wire_constant;
    -- flow-through select operator MUX_1407_inst
    MUX_1407_wire <= konst_1405_wire_constant when (read_from_4_1577(0) /=  '0') else konst_1406_wire_constant;
    -- flow-through select operator MUX_1455_inst
    MUX_1455_wire <= p1_valid_1421 when (EQ_u3_u1_1452_wire(0) /=  '0') else konst_1454_wire_constant;
    -- flow-through select operator MUX_1461_inst
    MUX_1461_wire <= p2_valid_1426 when (EQ_u3_u1_1458_wire(0) /=  '0') else konst_1460_wire_constant;
    -- flow-through select operator MUX_1468_inst
    MUX_1468_wire <= p3_valid_1431 when (EQ_u3_u1_1465_wire(0) /=  '0') else konst_1467_wire_constant;
    -- flow-through select operator MUX_1474_inst
    MUX_1474_wire <= p4_valid_1436 when (EQ_u3_u1_1471_wire(0) /=  '0') else konst_1473_wire_constant;
    -- flow-through select operator MUX_1505_inst
    MUX_1505_wire <= slice_1503_wire when (EQ_u3_u1_1501_wire(0) /=  '0') else konst_1504_wire_constant;
    -- flow-through select operator MUX_1512_inst
    MUX_1512_wire <= slice_1510_wire when (EQ_u3_u1_1508_wire(0) /=  '0') else konst_1511_wire_constant;
    -- flow-through select operator MUX_1520_inst
    MUX_1520_wire <= slice_1518_wire when (EQ_u3_u1_1516_wire(0) /=  '0') else konst_1519_wire_constant;
    -- flow-through select operator MUX_1527_inst
    MUX_1527_wire <= slice_1525_wire when (EQ_u3_u1_1523_wire(0) /=  '0') else konst_1526_wire_constant;
    -- flow-through select operator MUX_1531_inst
    next_active_packet_length_1532 <= OR_u8_u8_1529_wire when (started_new_packet_1496(0) /=  '0') else active_packet_length_1381;
    -- flow-through select operator MUX_1543_inst
    MUX_1543_wire <= SUB_u8_u8_1541_wire when (valid_active_pkt_word_read_1477(0) /=  '0') else down_counter_1353;
    -- flow-through select operator MUX_1544_inst
    next_down_counter_1545 <= SUB_u8_u8_1537_wire when (started_new_packet_1496(0) /=  '0') else MUX_1543_wire;
    -- flow-through select operator MUX_1585_inst
    MUX_1585_wire <= slice_1583_wire when (EQ_u3_u1_1581_wire(0) /=  '0') else konst_1584_wire_constant;
    -- flow-through select operator MUX_1592_inst
    MUX_1592_wire <= slice_1590_wire when (EQ_u3_u1_1588_wire(0) /=  '0') else konst_1591_wire_constant;
    -- flow-through select operator MUX_1600_inst
    MUX_1600_wire <= slice_1598_wire when (EQ_u3_u1_1596_wire(0) /=  '0') else konst_1599_wire_constant;
    -- flow-through select operator MUX_1607_inst
    MUX_1607_wire <= slice_1605_wire when (EQ_u3_u1_1603_wire(0) /=  '0') else konst_1606_wire_constant;
    -- flow-through select operator MUX_1617_inst
    MUX_1617_wire <= p1_valid_1421 when (EQ_u3_u1_1614_wire(0) /=  '0') else konst_1616_wire_constant;
    -- flow-through select operator MUX_1623_inst
    MUX_1623_wire <= p2_valid_1426 when (EQ_u3_u1_1620_wire(0) /=  '0') else konst_1622_wire_constant;
    -- flow-through select operator MUX_1630_inst
    MUX_1630_wire <= p3_valid_1431 when (EQ_u3_u1_1627_wire(0) /=  '0') else konst_1629_wire_constant;
    -- flow-through select operator MUX_1636_inst
    MUX_1636_wire <= p4_valid_1436 when (EQ_u3_u1_1633_wire(0) /=  '0') else konst_1635_wire_constant;
    -- flow-through slice operator slice_1503_inst
    slice_1503_wire <= pkt_1_e_word_1357(15 downto 8);
    -- flow-through slice operator slice_1510_inst
    slice_1510_wire <= pkt_2_e_word_1362(15 downto 8);
    -- flow-through slice operator slice_1518_inst
    slice_1518_wire <= pkt_3_e_word_1367(15 downto 8);
    -- flow-through slice operator slice_1525_inst
    slice_1525_wire <= pkt_4_e_word_1372(15 downto 8);
    -- flow-through slice operator slice_1583_inst
    slice_1583_wire <= pkt_1_e_word_1357(31 downto 0);
    -- flow-through slice operator slice_1590_inst
    slice_1590_wire <= pkt_2_e_word_1362(31 downto 0);
    -- flow-through slice operator slice_1598_inst
    slice_1598_wire <= pkt_3_e_word_1367(31 downto 0);
    -- flow-through slice operator slice_1605_inst
    slice_1605_wire <= pkt_4_e_word_1372(31 downto 0);
    next_active_packet_1487_1380_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_active_packet_1487_1380_buf_req_0;
      next_active_packet_1487_1380_buf_ack_0<= wack(0);
      rreq(0) <= next_active_packet_1487_1380_buf_req_1;
      next_active_packet_1487_1380_buf_ack_1<= rack(0);
      next_active_packet_1487_1380_buf : InterlockBuffer generic map ( -- 
        name => "next_active_packet_1487_1380_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_active_packet_1487,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_active_packet_1487_1380_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_active_packet_length_1532_1384_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_active_packet_length_1532_1384_buf_req_0;
      next_active_packet_length_1532_1384_buf_ack_0<= wack(0);
      rreq(0) <= next_active_packet_length_1532_1384_buf_req_1;
      next_active_packet_length_1532_1384_buf_ack_1<= rack(0);
      next_active_packet_length_1532_1384_buf : InterlockBuffer generic map ( -- 
        name => "next_active_packet_length_1532_1384_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_active_packet_length_1532,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_active_packet_length_1532_1384_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_down_counter_1545_1356_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_down_counter_1545_1356_buf_req_0;
      next_down_counter_1545_1356_buf_ack_0<= wack(0);
      rreq(0) <= next_down_counter_1545_1356_buf_req_1;
      next_down_counter_1545_1356_buf_ack_1<= rack(0);
      next_down_counter_1545_1356_buf : InterlockBuffer generic map ( -- 
        name => "next_down_counter_1545_1356_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_down_counter_1545,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_down_counter_1545_1356_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_priority_index_1487_1388_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_priority_index_1487_1388_buf_req_0;
      next_priority_index_1487_1388_buf_ack_0<= wack(0);
      rreq(0) <= next_priority_index_1487_1388_buf_req_1;
      next_priority_index_1487_1388_buf_ack_1<= rack(0);
      next_priority_index_1487_1388_buf : InterlockBuffer generic map ( -- 
        name => "next_priority_index_1487_1388_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 2,
        out_data_width => 2,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_priority_index_1487,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_priority_index_1487_1388_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1351_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1654_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1351_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1351_branch_req_0,
          ack0 => do_while_stmt_1351_branch_ack_0,
          ack1 => do_while_stmt_1351_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- flow through binary operator AND_u1_u1_1495_inst
    started_new_packet_1496 <= (NEQ_u3_u1_1491_wire and EQ_u8_u1_1494_wire);
    -- flow through binary operator BITSEL_u33_u1_1420_inst
    process(pkt_1_e_word_1357) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_1_e_word_1357, konst_1419_wire_constant, tmp_var);
      p1_valid_1421 <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u33_u1_1425_inst
    process(pkt_2_e_word_1362) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_2_e_word_1362, konst_1424_wire_constant, tmp_var);
      p2_valid_1426 <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u33_u1_1430_inst
    process(pkt_3_e_word_1367) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_3_e_word_1367, konst_1429_wire_constant, tmp_var);
      p3_valid_1431 <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u33_u1_1435_inst
    process(pkt_4_e_word_1372) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_4_e_word_1372, konst_1434_wire_constant, tmp_var);
      p4_valid_1436 <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1452_inst
    process(active_packet_1377) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1377, konst_1451_wire_constant, tmp_var);
      EQ_u3_u1_1452_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1458_inst
    process(active_packet_1377) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1377, konst_1457_wire_constant, tmp_var);
      EQ_u3_u1_1458_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1465_inst
    process(active_packet_1377) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1377, konst_1464_wire_constant, tmp_var);
      EQ_u3_u1_1465_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1471_inst
    process(active_packet_1377) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1377, konst_1470_wire_constant, tmp_var);
      EQ_u3_u1_1471_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1501_inst
    process(next_active_packet_1487) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1487, konst_1500_wire_constant, tmp_var);
      EQ_u3_u1_1501_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1508_inst
    process(next_active_packet_1487) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1487, konst_1507_wire_constant, tmp_var);
      EQ_u3_u1_1508_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1516_inst
    process(next_active_packet_1487) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1487, konst_1515_wire_constant, tmp_var);
      EQ_u3_u1_1516_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1523_inst
    process(next_active_packet_1487) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1487, konst_1522_wire_constant, tmp_var);
      EQ_u3_u1_1523_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1551_inst
    process(next_active_packet_1487) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1487, konst_1550_wire_constant, tmp_var);
      EQ_u3_u1_1551_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1559_inst
    process(next_active_packet_1487) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1487, konst_1558_wire_constant, tmp_var);
      EQ_u3_u1_1559_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1567_inst
    process(next_active_packet_1487) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1487, konst_1566_wire_constant, tmp_var);
      EQ_u3_u1_1567_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1575_inst
    process(next_active_packet_1487) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1487, konst_1574_wire_constant, tmp_var);
      EQ_u3_u1_1575_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1581_inst
    process(next_active_packet_1487) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1487, konst_1580_wire_constant, tmp_var);
      EQ_u3_u1_1581_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1588_inst
    process(next_active_packet_1487) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1487, konst_1587_wire_constant, tmp_var);
      EQ_u3_u1_1588_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1596_inst
    process(next_active_packet_1487) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1487, konst_1595_wire_constant, tmp_var);
      EQ_u3_u1_1596_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1603_inst
    process(next_active_packet_1487) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1487, konst_1602_wire_constant, tmp_var);
      EQ_u3_u1_1603_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1614_inst
    process(next_active_packet_1487) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1487, konst_1613_wire_constant, tmp_var);
      EQ_u3_u1_1614_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1620_inst
    process(next_active_packet_1487) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1487, konst_1619_wire_constant, tmp_var);
      EQ_u3_u1_1620_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1627_inst
    process(next_active_packet_1487) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1487, konst_1626_wire_constant, tmp_var);
      EQ_u3_u1_1627_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1633_inst
    process(next_active_packet_1487) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1487, konst_1632_wire_constant, tmp_var);
      EQ_u3_u1_1633_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u8_u1_1494_inst
    process(down_counter_1353) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(down_counter_1353, konst_1493_wire_constant, tmp_var);
      EQ_u8_u1_1494_wire <= tmp_var; --
    end process;
    -- flow through binary operator NEQ_u3_u1_1491_inst
    process(next_active_packet_1487) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(next_active_packet_1487, konst_1490_wire_constant, tmp_var);
      NEQ_u3_u1_1491_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1548_inst
    process(p1_valid_1421) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p1_valid_1421, tmp_var);
      NOT_u1_u1_1548_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1556_inst
    process(p2_valid_1426) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p2_valid_1426, tmp_var);
      NOT_u1_u1_1556_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1564_inst
    process(p3_valid_1431) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p3_valid_1431, tmp_var);
      NOT_u1_u1_1564_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1572_inst
    process(p4_valid_1436) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p4_valid_1436, tmp_var);
      NOT_u1_u1_1572_wire <= tmp_var; -- 
    end process;
    -- flow through binary operator OR_u1_u1_1462_inst
    OR_u1_u1_1462_wire <= (MUX_1455_wire or MUX_1461_wire);
    -- flow through binary operator OR_u1_u1_1475_inst
    OR_u1_u1_1475_wire <= (MUX_1468_wire or MUX_1474_wire);
    -- flow through binary operator OR_u1_u1_1476_inst
    valid_active_pkt_word_read_1477 <= (OR_u1_u1_1462_wire or OR_u1_u1_1475_wire);
    -- flow through binary operator OR_u1_u1_1552_inst
    read_from_1_1553 <= (NOT_u1_u1_1548_wire or EQ_u3_u1_1551_wire);
    -- flow through binary operator OR_u1_u1_1560_inst
    read_from_2_1561 <= (NOT_u1_u1_1556_wire or EQ_u3_u1_1559_wire);
    -- flow through binary operator OR_u1_u1_1568_inst
    read_from_3_1569 <= (NOT_u1_u1_1564_wire or EQ_u3_u1_1567_wire);
    -- flow through binary operator OR_u1_u1_1576_inst
    read_from_4_1577 <= (NOT_u1_u1_1572_wire or EQ_u3_u1_1575_wire);
    -- flow through binary operator OR_u1_u1_1624_inst
    OR_u1_u1_1624_wire <= (MUX_1617_wire or MUX_1623_wire);
    -- flow through binary operator OR_u1_u1_1637_inst
    OR_u1_u1_1637_wire <= (MUX_1630_wire or MUX_1636_wire);
    -- flow through binary operator OR_u1_u1_1638_inst
    send_flag_1639 <= (OR_u1_u1_1624_wire or OR_u1_u1_1637_wire);
    -- flow through binary operator OR_u32_u32_1593_inst
    OR_u32_u32_1593_wire <= (MUX_1585_wire or MUX_1592_wire);
    -- flow through binary operator OR_u32_u32_1608_inst
    OR_u32_u32_1608_wire <= (MUX_1600_wire or MUX_1607_wire);
    -- flow through binary operator OR_u32_u32_1609_inst
    data_to_out_1610 <= (OR_u32_u32_1593_wire or OR_u32_u32_1608_wire);
    -- flow through binary operator OR_u8_u8_1399_inst
    OR_u8_u8_1399_wire <= (MUX_1394_wire or MUX_1398_wire);
    -- flow through binary operator OR_u8_u8_1408_inst
    OR_u8_u8_1408_wire <= (MUX_1403_wire or MUX_1407_wire);
    -- flow through binary operator OR_u8_u8_1409_inst
    senderPort_1410 <= (OR_u8_u8_1399_wire or OR_u8_u8_1408_wire);
    -- flow through binary operator OR_u8_u8_1513_inst
    OR_u8_u8_1513_wire <= (MUX_1505_wire or MUX_1512_wire);
    -- flow through binary operator OR_u8_u8_1528_inst
    OR_u8_u8_1528_wire <= (MUX_1520_wire or MUX_1527_wire);
    -- flow through binary operator OR_u8_u8_1529_inst
    OR_u8_u8_1529_wire <= (OR_u8_u8_1513_wire or OR_u8_u8_1528_wire);
    -- flow through binary operator SUB_u8_u8_1537_inst
    SUB_u8_u8_1537_wire <= std_logic_vector(unsigned(next_active_packet_length_1532) - unsigned(konst_1536_wire_constant));
    -- flow through binary operator SUB_u8_u8_1541_inst
    SUB_u8_u8_1541_wire <= std_logic_vector(unsigned(down_counter_1353) - unsigned(konst_1540_wire_constant));
    -- shared inport operator group (0) : RPIPE_noblock_obuf_1_2_1361_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_1_2_1361_inst_req_0;
      RPIPE_noblock_obuf_1_2_1361_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_1_2_1361_inst_req_1;
      RPIPE_noblock_obuf_1_2_1361_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_1_1553(0);
      RPIPE_noblock_obuf_1_2_1361_wire <= data_out(32 downto 0);
      noblock_obuf_1_2_read_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_2_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_2_read_0: InputPortRevised -- 
        generic map ( name => "noblock_obuf_1_2_read_0", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_1_2_pipe_read_req(0),
          oack => noblock_obuf_1_2_pipe_read_ack(0),
          odata => noblock_obuf_1_2_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_noblock_obuf_2_2_1366_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_2_2_1366_inst_req_0;
      RPIPE_noblock_obuf_2_2_1366_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_2_2_1366_inst_req_1;
      RPIPE_noblock_obuf_2_2_1366_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_2_1561(0);
      RPIPE_noblock_obuf_2_2_1366_wire <= data_out(32 downto 0);
      noblock_obuf_2_2_read_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_2_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_2_read_1: InputPortRevised -- 
        generic map ( name => "noblock_obuf_2_2_read_1", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_2_2_pipe_read_req(0),
          oack => noblock_obuf_2_2_pipe_read_ack(0),
          odata => noblock_obuf_2_2_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_noblock_obuf_3_2_1371_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_3_2_1371_inst_req_0;
      RPIPE_noblock_obuf_3_2_1371_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_3_2_1371_inst_req_1;
      RPIPE_noblock_obuf_3_2_1371_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_3_1569(0);
      RPIPE_noblock_obuf_3_2_1371_wire <= data_out(32 downto 0);
      noblock_obuf_3_2_read_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_2_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_2_read_2: InputPortRevised -- 
        generic map ( name => "noblock_obuf_3_2_read_2", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_3_2_pipe_read_req(0),
          oack => noblock_obuf_3_2_pipe_read_ack(0),
          odata => noblock_obuf_3_2_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_noblock_obuf_4_2_1376_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_4_2_1376_inst_req_0;
      RPIPE_noblock_obuf_4_2_1376_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_4_2_1376_inst_req_1;
      RPIPE_noblock_obuf_4_2_1376_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_4_1577(0);
      RPIPE_noblock_obuf_4_2_1376_wire <= data_out(32 downto 0);
      noblock_obuf_4_2_read_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_2_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_2_read_3: InputPortRevised -- 
        generic map ( name => "noblock_obuf_4_2_read_3", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_4_2_pipe_read_req(0),
          oack => noblock_obuf_4_2_pipe_read_ack(0),
          odata => noblock_obuf_4_2_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_out_data_2_1641_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_out_data_2_1641_inst_req_0;
      WPIPE_out_data_2_1641_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_out_data_2_1641_inst_req_1;
      WPIPE_out_data_2_1641_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_flag_1639(0);
      data_in <= data_to_out_1610;
      out_data_2_write_0_gI: SplitGuardInterface generic map(name => "out_data_2_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      out_data_2_write_0: OutputPortRevised -- 
        generic map ( name => "out_data_2", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => out_data_2_pipe_write_req(0),
          oack => out_data_2_pipe_write_ack(0),
          odata => out_data_2_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_1416_call 
    updateCounter_call_group_0: Block -- 
      signal data_in: std_logic_vector(16 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1416_call_req_0;
      call_stmt_1416_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1416_call_req_1;
      call_stmt_1416_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      updateCounter_call_group_0_gI: SplitGuardInterface generic map(name => "updateCounter_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= senderPort_1410 & konst_1412_wire_constant & type_cast_1414_wire_constant;
      continue_1416 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 17,
        owidth => 17,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => updateCounter_call_reqs(0),
          ackR => updateCounter_call_acks(0),
          dataR => updateCounter_call_data(16 downto 0),
          tagR => updateCounter_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => updateCounter_return_acks(0), -- cross-over
          ackL => updateCounter_return_reqs(0), -- cross-over
          dataL => updateCounter_return_data(0 downto 0),
          tagL => updateCounter_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    volatile_operator_prioritySelect_4960: prioritySelect_Volatile port map(down_counter => down_counter_1353, active_packet => active_packet_1377, priority_index => priority_index_1385, p1_valid => p1_valid_1421, p2_valid => p2_valid_1426, p3_valid => p3_valid_1431, p4_valid => p4_valid_1436, next_active_packet => next_active_packet_1487, next_priority_index => next_priority_index_1487); 
    -- 
  end Block; -- data_path
  -- 
end outputPort_2_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity outputPort_3_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    noblock_obuf_1_3_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_3_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_3_3_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_3_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_4_3_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_3_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_2_3_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_3_pipe_read_data : in   std_logic_vector(32 downto 0);
    out_data_3_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_data_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_data_3_pipe_write_data : out  std_logic_vector(31 downto 0);
    updateCounter_call_reqs : out  std_logic_vector(0 downto 0);
    updateCounter_call_acks : in   std_logic_vector(0 downto 0);
    updateCounter_call_data : out  std_logic_vector(16 downto 0);
    updateCounter_call_tag  :  out  std_logic_vector(0 downto 0);
    updateCounter_return_reqs : out  std_logic_vector(0 downto 0);
    updateCounter_return_acks : in   std_logic_vector(0 downto 0);
    updateCounter_return_data : in   std_logic_vector(0 downto 0);
    updateCounter_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity outputPort_3_Daemon;
architecture outputPort_3_Daemon_arch of outputPort_3_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal outputPort_3_Daemon_CP_3266_start: Boolean;
  signal outputPort_3_Daemon_CP_3266_symbol: Boolean;
  -- volatile/operator module components. 
  component updateCounter is -- 
    generic (tag_length : integer); 
    port ( -- 
      input_port : in  std_logic_vector(7 downto 0);
      output_port : in  std_logic_vector(7 downto 0);
      up : in  std_logic_vector(0 downto 0);
      continue : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(3 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(1 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(1 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component prioritySelect_Volatile is -- 
    port ( -- 
      down_counter : in  std_logic_vector(7 downto 0);
      active_packet : in  std_logic_vector(2 downto 0);
      priority_index : in  std_logic_vector(1 downto 0);
      p1_valid : in  std_logic_vector(0 downto 0);
      p2_valid : in  std_logic_vector(0 downto 0);
      p3_valid : in  std_logic_vector(0 downto 0);
      p4_valid : in  std_logic_vector(0 downto 0);
      next_active_packet : out  std_logic_vector(2 downto 0);
      next_priority_index : out  std_logic_vector(1 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal phi_stmt_1680_req_0 : boolean;
  signal next_down_counter_1853_1664_buf_req_1 : boolean;
  signal RPIPE_noblock_obuf_1_3_1669_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_3_3_1679_inst_ack_1 : boolean;
  signal RPIPE_noblock_obuf_3_3_1679_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_3_3_1679_inst_req_1 : boolean;
  signal next_down_counter_1853_1664_buf_ack_1 : boolean;
  signal RPIPE_noblock_obuf_3_3_1679_inst_ack_0 : boolean;
  signal phi_stmt_1661_req_0 : boolean;
  signal phi_stmt_1665_req_1 : boolean;
  signal RPIPE_noblock_obuf_2_3_1674_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_2_3_1674_inst_ack_0 : boolean;
  signal phi_stmt_1665_req_0 : boolean;
  signal phi_stmt_1665_ack_0 : boolean;
  signal phi_stmt_1670_req_1 : boolean;
  signal phi_stmt_1675_ack_0 : boolean;
  signal RPIPE_noblock_obuf_2_3_1674_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_2_3_1674_inst_ack_1 : boolean;
  signal phi_stmt_1661_req_1 : boolean;
  signal phi_stmt_1670_req_0 : boolean;
  signal phi_stmt_1675_req_1 : boolean;
  signal RPIPE_noblock_obuf_1_3_1669_inst_ack_1 : boolean;
  signal do_while_stmt_1659_branch_req_0 : boolean;
  signal RPIPE_noblock_obuf_1_3_1669_inst_req_0 : boolean;
  signal phi_stmt_1675_req_0 : boolean;
  signal RPIPE_noblock_obuf_1_3_1669_inst_ack_0 : boolean;
  signal phi_stmt_1680_ack_0 : boolean;
  signal phi_stmt_1685_req_1 : boolean;
  signal next_down_counter_1853_1664_buf_ack_0 : boolean;
  signal next_down_counter_1853_1664_buf_req_0 : boolean;
  signal RPIPE_noblock_obuf_4_3_1684_inst_req_0 : boolean;
  signal phi_stmt_1685_ack_0 : boolean;
  signal next_active_packet_1795_1688_buf_req_1 : boolean;
  signal next_active_packet_1795_1688_buf_ack_1 : boolean;
  signal next_active_packet_1795_1688_buf_ack_0 : boolean;
  signal next_active_packet_1795_1688_buf_req_0 : boolean;
  signal RPIPE_noblock_obuf_4_3_1684_inst_ack_1 : boolean;
  signal phi_stmt_1680_req_1 : boolean;
  signal phi_stmt_1685_req_0 : boolean;
  signal RPIPE_noblock_obuf_4_3_1684_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_4_3_1684_inst_ack_0 : boolean;
  signal phi_stmt_1670_ack_0 : boolean;
  signal phi_stmt_1661_ack_0 : boolean;
  signal phi_stmt_1689_req_1 : boolean;
  signal phi_stmt_1689_req_0 : boolean;
  signal phi_stmt_1689_ack_0 : boolean;
  signal next_active_packet_length_1840_1692_buf_req_0 : boolean;
  signal next_active_packet_length_1840_1692_buf_ack_0 : boolean;
  signal next_active_packet_length_1840_1692_buf_req_1 : boolean;
  signal next_active_packet_length_1840_1692_buf_ack_1 : boolean;
  signal phi_stmt_1693_req_0 : boolean;
  signal phi_stmt_1693_req_1 : boolean;
  signal phi_stmt_1693_ack_0 : boolean;
  signal next_priority_index_1795_1695_buf_req_0 : boolean;
  signal next_priority_index_1795_1695_buf_ack_0 : boolean;
  signal next_priority_index_1795_1695_buf_req_1 : boolean;
  signal next_priority_index_1795_1695_buf_ack_1 : boolean;
  signal call_stmt_1724_call_req_0 : boolean;
  signal call_stmt_1724_call_ack_0 : boolean;
  signal call_stmt_1724_call_req_1 : boolean;
  signal call_stmt_1724_call_ack_1 : boolean;
  signal WPIPE_out_data_3_1949_inst_req_0 : boolean;
  signal WPIPE_out_data_3_1949_inst_ack_0 : boolean;
  signal WPIPE_out_data_3_1949_inst_req_1 : boolean;
  signal WPIPE_out_data_3_1949_inst_ack_1 : boolean;
  signal do_while_stmt_1659_branch_ack_0 : boolean;
  signal do_while_stmt_1659_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "outputPort_3_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  outputPort_3_Daemon_CP_3266_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "outputPort_3_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_3_Daemon_CP_3266_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= outputPort_3_Daemon_CP_3266_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_3_Daemon_CP_3266_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  outputPort_3_Daemon_CP_3266: Block -- control-path 
    signal outputPort_3_Daemon_CP_3266_elements: BooleanArray(185 downto 0);
    -- 
  begin -- 
    outputPort_3_Daemon_CP_3266_elements(0) <= outputPort_3_Daemon_CP_3266_start;
    outputPort_3_Daemon_CP_3266_symbol <= outputPort_3_Daemon_CP_3266_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1658/branch_block_stmt_1658__entry__
      -- CP-element group 0: 	 branch_block_stmt_1658/$entry
      -- CP-element group 0: 	 branch_block_stmt_1658/do_while_stmt_1659__entry__
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	185 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_1658/do_while_stmt_1659__exit__
      -- CP-element group 1: 	 branch_block_stmt_1658/branch_block_stmt_1658__exit__
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1658/$exit
      -- 
    outputPort_3_Daemon_CP_3266_elements(1) <= outputPort_3_Daemon_CP_3266_elements(185);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659__entry__
      -- CP-element group 2: 	 branch_block_stmt_1658/do_while_stmt_1659/$entry
      -- 
    outputPort_3_Daemon_CP_3266_elements(2) <= outputPort_3_Daemon_CP_3266_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	185 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659__exit__
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1658/do_while_stmt_1659/loop_back
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	184 
    -- CP-element group 5: 	183 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1658/do_while_stmt_1659/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1658/do_while_stmt_1659/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1658/do_while_stmt_1659/loop_taken/$entry
      -- 
    outputPort_3_Daemon_CP_3266_elements(5) <= outputPort_3_Daemon_CP_3266_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	182 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1658/do_while_stmt_1659/loop_body_done
      -- 
    outputPort_3_Daemon_CP_3266_elements(6) <= outputPort_3_Daemon_CP_3266_elements(182);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	124 
    -- CP-element group 7: 	161 
    -- CP-element group 7: 	104 
    -- CP-element group 7: 	83 
    -- CP-element group 7: 	22 
    -- CP-element group 7: 	41 
    -- CP-element group 7: 	143 
    -- CP-element group 7: 	62 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/back_edge_to_loop_body
      -- 
    outputPort_3_Daemon_CP_3266_elements(7) <= outputPort_3_Daemon_CP_3266_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	126 
    -- CP-element group 8: 	163 
    -- CP-element group 8: 	106 
    -- CP-element group 8: 	85 
    -- CP-element group 8: 	24 
    -- CP-element group 8: 	43 
    -- CP-element group 8: 	145 
    -- CP-element group 8: 	64 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/first_time_through_loop_body
      -- 
    outputPort_3_Daemon_CP_3266_elements(8) <= outputPort_3_Daemon_CP_3266_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	156 
    -- CP-element group 9: 	157 
    -- CP-element group 9: 	137 
    -- CP-element group 9: 	138 
    -- CP-element group 9: 	119 
    -- CP-element group 9: 	120 
    -- CP-element group 9: 	181 
    -- CP-element group 9: 	77 
    -- CP-element group 9: 	78 
    -- CP-element group 9: 	98 
    -- CP-element group 9: 	99 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	17 
    -- CP-element group 9: 	35 
    -- CP-element group 9: 	36 
    -- CP-element group 9: 	56 
    -- CP-element group 9: 	57 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/loop_body_start
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	181 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/condition_evaluated
      -- 
    condition_evaluated_3290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(10), ack => do_while_stmt_1659_branch_req_0); -- 
    outputPort_3_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(181) & outputPort_3_Daemon_CP_3266_elements(15);
      gj_outputPort_3_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	156 
    -- CP-element group 11: 	137 
    -- CP-element group 11: 	119 
    -- CP-element group 11: 	77 
    -- CP-element group 11: 	98 
    -- CP-element group 11: 	16 
    -- CP-element group 11: 	35 
    -- CP-element group 11: 	56 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	121 
    -- CP-element group 11: 	139 
    -- CP-element group 11: 	100 
    -- CP-element group 11: 	79 
    -- CP-element group 11: 	18 
    -- CP-element group 11: 	37 
    -- CP-element group 11: 	58 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1693_sample_start__ps
      -- CP-element group 11: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/aggregated_phi_sample_req
      -- 
    outputPort_3_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 1);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(156) & outputPort_3_Daemon_CP_3266_elements(137) & outputPort_3_Daemon_CP_3266_elements(119) & outputPort_3_Daemon_CP_3266_elements(77) & outputPort_3_Daemon_CP_3266_elements(98) & outputPort_3_Daemon_CP_3266_elements(16) & outputPort_3_Daemon_CP_3266_elements(35) & outputPort_3_Daemon_CP_3266_elements(56) & outputPort_3_Daemon_CP_3266_elements(15);
      gj_outputPort_3_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	122 
    -- CP-element group 12: 	158 
    -- CP-element group 12: 	140 
    -- CP-element group 12: 	101 
    -- CP-element group 12: 	80 
    -- CP-element group 12: 	19 
    -- CP-element group 12: 	38 
    -- CP-element group 12: 	59 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	182 
    -- CP-element group 12: 	13 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	156 
    -- CP-element group 12: 	137 
    -- CP-element group 12: 	119 
    -- CP-element group 12: 	77 
    -- CP-element group 12: 	98 
    -- CP-element group 12: 	16 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	56 
    -- CP-element group 12:  members (9) 
      -- CP-element group 12: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1680_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1675_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1665_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1670_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1661_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1685_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1689_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1693_sample_completed_
      -- 
    outputPort_3_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(122) & outputPort_3_Daemon_CP_3266_elements(158) & outputPort_3_Daemon_CP_3266_elements(140) & outputPort_3_Daemon_CP_3266_elements(101) & outputPort_3_Daemon_CP_3266_elements(80) & outputPort_3_Daemon_CP_3266_elements(19) & outputPort_3_Daemon_CP_3266_elements(38) & outputPort_3_Daemon_CP_3266_elements(59);
      gj_outputPort_3_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	182 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/aggregated_phi_sample_ack_d
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(13) is a control-delay.
    cp_element_13_delay: control_delay_element  generic map(name => " 13_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_3266_elements(12), ack => outputPort_3_Daemon_CP_3266_elements(13), clk => clk, reset =>reset);
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	157 
    -- CP-element group 14: 	138 
    -- CP-element group 14: 	120 
    -- CP-element group 14: 	78 
    -- CP-element group 14: 	99 
    -- CP-element group 14: 	17 
    -- CP-element group 14: 	36 
    -- CP-element group 14: 	57 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	159 
    -- CP-element group 14: 	141 
    -- CP-element group 14: 	102 
    -- CP-element group 14: 	81 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	39 
    -- CP-element group 14: 	60 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/aggregated_phi_update_req
      -- CP-element group 14: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1685_update_start__ps
      -- 
    outputPort_3_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(157) & outputPort_3_Daemon_CP_3266_elements(138) & outputPort_3_Daemon_CP_3266_elements(120) & outputPort_3_Daemon_CP_3266_elements(78) & outputPort_3_Daemon_CP_3266_elements(99) & outputPort_3_Daemon_CP_3266_elements(17) & outputPort_3_Daemon_CP_3266_elements(36) & outputPort_3_Daemon_CP_3266_elements(57);
      gj_outputPort_3_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	123 
    -- CP-element group 15: 	160 
    -- CP-element group 15: 	142 
    -- CP-element group 15: 	82 
    -- CP-element group 15: 	103 
    -- CP-element group 15: 	21 
    -- CP-element group 15: 	40 
    -- CP-element group 15: 	61 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/aggregated_phi_update_ack
      -- 
    outputPort_3_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 7);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(123) & outputPort_3_Daemon_CP_3266_elements(160) & outputPort_3_Daemon_CP_3266_elements(142) & outputPort_3_Daemon_CP_3266_elements(82) & outputPort_3_Daemon_CP_3266_elements(103) & outputPort_3_Daemon_CP_3266_elements(21) & outputPort_3_Daemon_CP_3266_elements(40) & outputPort_3_Daemon_CP_3266_elements(61);
      gj_outputPort_3_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	11 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1661_sample_start_
      -- 
    outputPort_3_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(9) & outputPort_3_Daemon_CP_3266_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	9 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	176 
    -- CP-element group 17: 	179 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	14 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1661_update_start_
      -- 
    outputPort_3_Daemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(9) & outputPort_3_Daemon_CP_3266_elements(176) & outputPort_3_Daemon_CP_3266_elements(179);
      gj_outputPort_3_Daemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	11 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1661_sample_start__ps
      -- 
    outputPort_3_Daemon_CP_3266_elements(18) <= outputPort_3_Daemon_CP_3266_elements(11);
    -- CP-element group 19:  join  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	12 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1661_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(19) is bound as output of CP function.
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	14 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1661_update_start__ps
      -- 
    outputPort_3_Daemon_CP_3266_elements(20) <= outputPort_3_Daemon_CP_3266_elements(14);
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	174 
    -- CP-element group 21: 	178 
    -- CP-element group 21: 	15 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1661_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1661_update_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(21) is bound as output of CP function.
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	7 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1661_loopback_trigger
      -- 
    outputPort_3_Daemon_CP_3266_elements(22) <= outputPort_3_Daemon_CP_3266_elements(7);
    -- CP-element group 23:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1661_loopback_sample_req
      -- CP-element group 23: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1661_loopback_sample_req_ps
      -- 
    phi_stmt_1661_loopback_sample_req_3306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1661_loopback_sample_req_3306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(23), ack => phi_stmt_1661_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(23) is bound as output of CP function.
    -- CP-element group 24:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	8 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1661_entry_trigger
      -- 
    outputPort_3_Daemon_CP_3266_elements(24) <= outputPort_3_Daemon_CP_3266_elements(8);
    -- CP-element group 25:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1661_entry_sample_req_ps
      -- CP-element group 25: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1661_entry_sample_req
      -- 
    phi_stmt_1661_entry_sample_req_3309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1661_entry_sample_req_3309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(25), ack => phi_stmt_1661_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1661_phi_mux_ack_ps
      -- CP-element group 26: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1661_phi_mux_ack
      -- 
    phi_stmt_1661_phi_mux_ack_3312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1661_ack_0, ack => outputPort_3_Daemon_CP_3266_elements(26)); -- 
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_8_1663_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_8_1663_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_8_1663_sample_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_8_1663_sample_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_8_1663_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_8_1663_update_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	30 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_8_1663_update_completed__ps
      -- 
    outputPort_3_Daemon_CP_3266_elements(29) <= outputPort_3_Daemon_CP_3266_elements(30);
    -- CP-element group 30:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	29 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_8_1663_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(30) is a control-delay.
    cp_element_30_delay: control_delay_element  generic map(name => " 30_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_3266_elements(28), ack => outputPort_3_Daemon_CP_3266_elements(30), clk => clk, reset =>reset);
    -- CP-element group 31:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_down_counter_1664_Sample/req
      -- CP-element group 31: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_down_counter_1664_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_down_counter_1664_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_down_counter_1664_sample_start__ps
      -- 
    req_3333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(31), ack => next_down_counter_1853_1664_buf_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_down_counter_1664_Update/req
      -- CP-element group 32: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_down_counter_1664_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_down_counter_1664_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_down_counter_1664_update_start__ps
      -- 
    req_3338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(32), ack => next_down_counter_1853_1664_buf_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_down_counter_1664_Sample/ack
      -- CP-element group 33: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_down_counter_1664_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_down_counter_1664_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_down_counter_1664_sample_completed__ps
      -- 
    ack_3334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_1853_1664_buf_ack_0, ack => outputPort_3_Daemon_CP_3266_elements(33)); -- 
    -- CP-element group 34:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_down_counter_1664_Update/ack
      -- CP-element group 34: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_down_counter_1664_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_down_counter_1664_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_down_counter_1664_update_completed__ps
      -- 
    ack_3339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_1853_1664_buf_ack_1, ack => outputPort_3_Daemon_CP_3266_elements(34)); -- 
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	12 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	11 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1665_sample_start_
      -- 
    outputPort_3_Daemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(9) & outputPort_3_Daemon_CP_3266_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	9 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	176 
    -- CP-element group 36: 	179 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	14 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1665_update_start_
      -- 
    outputPort_3_Daemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(9) & outputPort_3_Daemon_CP_3266_elements(176) & outputPort_3_Daemon_CP_3266_elements(179);
      gj_outputPort_3_Daemon_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	11 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1665_sample_start__ps
      -- 
    outputPort_3_Daemon_CP_3266_elements(37) <= outputPort_3_Daemon_CP_3266_elements(11);
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	12 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1665_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(38) is bound as output of CP function.
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	14 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1665_update_start__ps
      -- 
    outputPort_3_Daemon_CP_3266_elements(39) <= outputPort_3_Daemon_CP_3266_elements(14);
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	174 
    -- CP-element group 40: 	178 
    -- CP-element group 40: 	15 
    -- CP-element group 40:  members (2) 
      -- CP-element group 40: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1665_update_completed__ps
      -- CP-element group 40: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1665_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(40) is bound as output of CP function.
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	7 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1665_loopback_trigger
      -- 
    outputPort_3_Daemon_CP_3266_elements(41) <= outputPort_3_Daemon_CP_3266_elements(7);
    -- CP-element group 42:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1665_loopback_sample_req
      -- CP-element group 42: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1665_loopback_sample_req_ps
      -- 
    phi_stmt_1665_loopback_sample_req_3350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1665_loopback_sample_req_3350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(42), ack => phi_stmt_1665_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(42) is bound as output of CP function.
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	8 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1665_entry_trigger
      -- 
    outputPort_3_Daemon_CP_3266_elements(43) <= outputPort_3_Daemon_CP_3266_elements(8);
    -- CP-element group 44:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1665_entry_sample_req
      -- CP-element group 44: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1665_entry_sample_req_ps
      -- 
    phi_stmt_1665_entry_sample_req_3353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1665_entry_sample_req_3353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(44), ack => phi_stmt_1665_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(44) is bound as output of CP function.
    -- CP-element group 45:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1665_phi_mux_ack
      -- CP-element group 45: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1665_phi_mux_ack_ps
      -- 
    phi_stmt_1665_phi_mux_ack_3356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1665_ack_0, ack => outputPort_3_Daemon_CP_3266_elements(45)); -- 
    -- CP-element group 46:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (4) 
      -- CP-element group 46: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1667_sample_start__ps
      -- CP-element group 46: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1667_sample_completed__ps
      -- CP-element group 46: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1667_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1667_sample_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1667_update_start__ps
      -- CP-element group 47: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1667_update_start_
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	49 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1667_update_completed__ps
      -- 
    outputPort_3_Daemon_CP_3266_elements(48) <= outputPort_3_Daemon_CP_3266_elements(49);
    -- CP-element group 49:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	48 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1667_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(49) is a control-delay.
    cp_element_49_delay: control_delay_element  generic map(name => " 49_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_3266_elements(47), ack => outputPort_3_Daemon_CP_3266_elements(49), clk => clk, reset =>reset);
    -- CP-element group 50:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_1_3_1669_sample_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_1_3_1669_update_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(51) is bound as output of CP function.
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	55 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_1_3_1669_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_1_3_1669_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_1_3_1669_Sample/rr
      -- 
    rr_3377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(52), ack => RPIPE_noblock_obuf_1_3_1669_inst_req_0); -- 
    outputPort_3_Daemon_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(50) & outputPort_3_Daemon_CP_3266_elements(55);
      gj_outputPort_3_Daemon_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: 	54 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_1_3_1669_Update/cr
      -- CP-element group 53: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_1_3_1669_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_1_3_1669_update_start_
      -- 
    cr_3382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(53), ack => RPIPE_noblock_obuf_1_3_1669_inst_req_1); -- 
    outputPort_3_Daemon_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(51) & outputPort_3_Daemon_CP_3266_elements(54);
      gj_outputPort_3_Daemon_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	53 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_1_3_1669_sample_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_1_3_1669_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_1_3_1669_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_1_3_1669_Sample/ra
      -- 
    ra_3378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_3_1669_inst_ack_0, ack => outputPort_3_Daemon_CP_3266_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: marked-successors 
    -- CP-element group 55: 	52 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_1_3_1669_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_1_3_1669_update_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_1_3_1669_Update/ca
      -- CP-element group 55: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_1_3_1669_update_completed_
      -- 
    ca_3383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_3_1669_inst_ack_1, ack => outputPort_3_Daemon_CP_3266_elements(55)); -- 
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	9 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	12 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	11 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1670_sample_start_
      -- 
    outputPort_3_Daemon_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(9) & outputPort_3_Daemon_CP_3266_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  join  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	9 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	176 
    -- CP-element group 57: 	179 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	14 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1670_update_start_
      -- 
    outputPort_3_Daemon_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(9) & outputPort_3_Daemon_CP_3266_elements(176) & outputPort_3_Daemon_CP_3266_elements(179);
      gj_outputPort_3_Daemon_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	11 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1670_sample_start__ps
      -- 
    outputPort_3_Daemon_CP_3266_elements(58) <= outputPort_3_Daemon_CP_3266_elements(11);
    -- CP-element group 59:  join  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	12 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1670_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(59) is bound as output of CP function.
    -- CP-element group 60:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	14 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1670_update_start__ps
      -- 
    outputPort_3_Daemon_CP_3266_elements(60) <= outputPort_3_Daemon_CP_3266_elements(14);
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	174 
    -- CP-element group 61: 	178 
    -- CP-element group 61: 	15 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1670_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1670_update_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(61) is bound as output of CP function.
    -- CP-element group 62:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	7 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1670_loopback_trigger
      -- 
    outputPort_3_Daemon_CP_3266_elements(62) <= outputPort_3_Daemon_CP_3266_elements(7);
    -- CP-element group 63:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1670_loopback_sample_req
      -- CP-element group 63: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1670_loopback_sample_req_ps
      -- 
    phi_stmt_1670_loopback_sample_req_3394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1670_loopback_sample_req_3394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(63), ack => phi_stmt_1670_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(63) is bound as output of CP function.
    -- CP-element group 64:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	8 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1670_entry_trigger
      -- 
    outputPort_3_Daemon_CP_3266_elements(64) <= outputPort_3_Daemon_CP_3266_elements(8);
    -- CP-element group 65:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1670_entry_sample_req
      -- CP-element group 65: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1670_entry_sample_req_ps
      -- 
    phi_stmt_1670_entry_sample_req_3397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1670_entry_sample_req_3397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(65), ack => phi_stmt_1670_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(65) is bound as output of CP function.
    -- CP-element group 66:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1670_phi_mux_ack_ps
      -- CP-element group 66: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1670_phi_mux_ack
      -- 
    phi_stmt_1670_phi_mux_ack_3400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1670_ack_0, ack => outputPort_3_Daemon_CP_3266_elements(66)); -- 
    -- CP-element group 67:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1672_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1672_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1672_sample_completed__ps
      -- CP-element group 67: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1672_sample_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1672_update_start_
      -- CP-element group 68: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1672_update_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	70 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1672_update_completed__ps
      -- 
    outputPort_3_Daemon_CP_3266_elements(69) <= outputPort_3_Daemon_CP_3266_elements(70);
    -- CP-element group 70:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	69 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1672_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(70) is a control-delay.
    cp_element_70_delay: control_delay_element  generic map(name => " 70_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_3266_elements(68), ack => outputPort_3_Daemon_CP_3266_elements(70), clk => clk, reset =>reset);
    -- CP-element group 71:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_2_3_1674_sample_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(71) is bound as output of CP function.
    -- CP-element group 72:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_2_3_1674_update_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(72) is bound as output of CP function.
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: marked-predecessors 
    -- CP-element group 73: 	76 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_2_3_1674_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_2_3_1674_Sample/rr
      -- CP-element group 73: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_2_3_1674_sample_start_
      -- 
    rr_3421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(73), ack => RPIPE_noblock_obuf_2_3_1674_inst_req_0); -- 
    outputPort_3_Daemon_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(71) & outputPort_3_Daemon_CP_3266_elements(76);
      gj_outputPort_3_Daemon_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: 	75 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_2_3_1674_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_2_3_1674_Update/cr
      -- CP-element group 74: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_2_3_1674_update_start_
      -- 
    cr_3426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(74), ack => RPIPE_noblock_obuf_2_3_1674_inst_req_1); -- 
    outputPort_3_Daemon_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(72) & outputPort_3_Daemon_CP_3266_elements(75);
      gj_outputPort_3_Daemon_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	74 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_2_3_1674_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_2_3_1674_Sample/ra
      -- CP-element group 75: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_2_3_1674_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_2_3_1674_sample_completed__ps
      -- 
    ra_3422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_3_1674_inst_ack_0, ack => outputPort_3_Daemon_CP_3266_elements(75)); -- 
    -- CP-element group 76:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: marked-successors 
    -- CP-element group 76: 	73 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_2_3_1674_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_2_3_1674_Update/ca
      -- CP-element group 76: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_2_3_1674_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_2_3_1674_update_completed__ps
      -- 
    ca_3427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_3_1674_inst_ack_1, ack => outputPort_3_Daemon_CP_3266_elements(76)); -- 
    -- CP-element group 77:  join  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	9 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	12 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	11 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1675_sample_start_
      -- 
    outputPort_3_Daemon_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(9) & outputPort_3_Daemon_CP_3266_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  join  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	9 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	176 
    -- CP-element group 78: 	179 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	14 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1675_update_start_
      -- 
    outputPort_3_Daemon_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(9) & outputPort_3_Daemon_CP_3266_elements(176) & outputPort_3_Daemon_CP_3266_elements(179);
      gj_outputPort_3_Daemon_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	11 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1675_sample_start__ps
      -- 
    outputPort_3_Daemon_CP_3266_elements(79) <= outputPort_3_Daemon_CP_3266_elements(11);
    -- CP-element group 80:  join  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	12 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1675_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(80) is bound as output of CP function.
    -- CP-element group 81:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	14 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1675_update_start__ps
      -- 
    outputPort_3_Daemon_CP_3266_elements(81) <= outputPort_3_Daemon_CP_3266_elements(14);
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	174 
    -- CP-element group 82: 	178 
    -- CP-element group 82: 	15 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1675_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1675_update_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(82) is bound as output of CP function.
    -- CP-element group 83:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	7 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1675_loopback_trigger
      -- 
    outputPort_3_Daemon_CP_3266_elements(83) <= outputPort_3_Daemon_CP_3266_elements(7);
    -- CP-element group 84:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1675_loopback_sample_req
      -- CP-element group 84: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1675_loopback_sample_req_ps
      -- 
    phi_stmt_1675_loopback_sample_req_3438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1675_loopback_sample_req_3438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(84), ack => phi_stmt_1675_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(84) is bound as output of CP function.
    -- CP-element group 85:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	8 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1675_entry_trigger
      -- 
    outputPort_3_Daemon_CP_3266_elements(85) <= outputPort_3_Daemon_CP_3266_elements(8);
    -- CP-element group 86:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1675_entry_sample_req_ps
      -- CP-element group 86: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1675_entry_sample_req
      -- 
    phi_stmt_1675_entry_sample_req_3441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1675_entry_sample_req_3441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(86), ack => phi_stmt_1675_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(86) is bound as output of CP function.
    -- CP-element group 87:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1675_phi_mux_ack
      -- CP-element group 87: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1675_phi_mux_ack_ps
      -- 
    phi_stmt_1675_phi_mux_ack_3444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1675_ack_0, ack => outputPort_3_Daemon_CP_3266_elements(87)); -- 
    -- CP-element group 88:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (4) 
      -- CP-element group 88: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1677_sample_start__ps
      -- CP-element group 88: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1677_sample_completed__ps
      -- CP-element group 88: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1677_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1677_sample_start_
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1677_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1677_update_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(89) is bound as output of CP function.
    -- CP-element group 90:  join  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	91 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1677_update_completed__ps
      -- 
    outputPort_3_Daemon_CP_3266_elements(90) <= outputPort_3_Daemon_CP_3266_elements(91);
    -- CP-element group 91:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	90 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1677_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(91) is a control-delay.
    cp_element_91_delay: control_delay_element  generic map(name => " 91_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_3266_elements(89), ack => outputPort_3_Daemon_CP_3266_elements(91), clk => clk, reset =>reset);
    -- CP-element group 92:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_3_3_1679_sample_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(92) is bound as output of CP function.
    -- CP-element group 93:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_3_3_1679_update_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(93) is bound as output of CP function.
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	97 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_3_3_1679_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_3_3_1679_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_3_3_1679_Sample/rr
      -- 
    rr_3465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(94), ack => RPIPE_noblock_obuf_3_3_1679_inst_req_0); -- 
    outputPort_3_Daemon_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(92) & outputPort_3_Daemon_CP_3266_elements(97);
      gj_outputPort_3_Daemon_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: 	96 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_3_3_1679_Update/cr
      -- CP-element group 95: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_3_3_1679_Update/$entry
      -- CP-element group 95: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_3_3_1679_update_start_
      -- 
    cr_3470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(95), ack => RPIPE_noblock_obuf_3_3_1679_inst_req_1); -- 
    outputPort_3_Daemon_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(93) & outputPort_3_Daemon_CP_3266_elements(96);
      gj_outputPort_3_Daemon_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	95 
    -- CP-element group 96:  members (4) 
      -- CP-element group 96: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_3_3_1679_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_3_3_1679_sample_completed__ps
      -- CP-element group 96: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_3_3_1679_Sample/ra
      -- CP-element group 96: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_3_3_1679_sample_completed_
      -- 
    ra_3466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_3_1679_inst_ack_0, ack => outputPort_3_Daemon_CP_3266_elements(96)); -- 
    -- CP-element group 97:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: marked-successors 
    -- CP-element group 97: 	94 
    -- CP-element group 97:  members (4) 
      -- CP-element group 97: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_3_3_1679_Update/ca
      -- CP-element group 97: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_3_3_1679_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_3_3_1679_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_3_3_1679_update_completed__ps
      -- 
    ca_3471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_3_1679_inst_ack_1, ack => outputPort_3_Daemon_CP_3266_elements(97)); -- 
    -- CP-element group 98:  join  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	9 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	12 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	11 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1680_sample_start_
      -- 
    outputPort_3_Daemon_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(9) & outputPort_3_Daemon_CP_3266_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  join  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	9 
    -- CP-element group 99: marked-predecessors 
    -- CP-element group 99: 	176 
    -- CP-element group 99: 	179 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	14 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1680_update_start_
      -- 
    outputPort_3_Daemon_cp_element_group_99: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_99"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(9) & outputPort_3_Daemon_CP_3266_elements(176) & outputPort_3_Daemon_CP_3266_elements(179);
      gj_outputPort_3_Daemon_cp_element_group_99 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(99), clk => clk, reset => reset); --
    end block;
    -- CP-element group 100:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	11 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1680_sample_start__ps
      -- 
    outputPort_3_Daemon_CP_3266_elements(100) <= outputPort_3_Daemon_CP_3266_elements(11);
    -- CP-element group 101:  join  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	12 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1680_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(101) is bound as output of CP function.
    -- CP-element group 102:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	14 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1680_update_start__ps
      -- 
    outputPort_3_Daemon_CP_3266_elements(102) <= outputPort_3_Daemon_CP_3266_elements(14);
    -- CP-element group 103:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	174 
    -- CP-element group 103: 	178 
    -- CP-element group 103: 	15 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1680_update_completed__ps
      -- CP-element group 103: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1680_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(103) is bound as output of CP function.
    -- CP-element group 104:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	7 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1680_loopback_trigger
      -- 
    outputPort_3_Daemon_CP_3266_elements(104) <= outputPort_3_Daemon_CP_3266_elements(7);
    -- CP-element group 105:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1680_loopback_sample_req_ps
      -- CP-element group 105: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1680_loopback_sample_req
      -- 
    phi_stmt_1680_loopback_sample_req_3482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1680_loopback_sample_req_3482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(105), ack => phi_stmt_1680_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(105) is bound as output of CP function.
    -- CP-element group 106:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	8 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1680_entry_trigger
      -- 
    outputPort_3_Daemon_CP_3266_elements(106) <= outputPort_3_Daemon_CP_3266_elements(8);
    -- CP-element group 107:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1680_entry_sample_req
      -- CP-element group 107: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1680_entry_sample_req_ps
      -- 
    phi_stmt_1680_entry_sample_req_3485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1680_entry_sample_req_3485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(107), ack => phi_stmt_1680_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(107) is bound as output of CP function.
    -- CP-element group 108:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1680_phi_mux_ack_ps
      -- CP-element group 108: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1680_phi_mux_ack
      -- 
    phi_stmt_1680_phi_mux_ack_3488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1680_ack_0, ack => outputPort_3_Daemon_CP_3266_elements(108)); -- 
    -- CP-element group 109:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (4) 
      -- CP-element group 109: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1682_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1682_sample_completed__ps
      -- CP-element group 109: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1682_sample_start__ps
      -- CP-element group 109: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1682_sample_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(109) is bound as output of CP function.
    -- CP-element group 110:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1682_update_start__ps
      -- CP-element group 110: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1682_update_start_
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(110) is bound as output of CP function.
    -- CP-element group 111:  join  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1682_update_completed__ps
      -- 
    outputPort_3_Daemon_CP_3266_elements(111) <= outputPort_3_Daemon_CP_3266_elements(112);
    -- CP-element group 112:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	111 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_33_1682_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(112) is a control-delay.
    cp_element_112_delay: control_delay_element  generic map(name => " 112_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_3266_elements(110), ack => outputPort_3_Daemon_CP_3266_elements(112), clk => clk, reset =>reset);
    -- CP-element group 113:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_4_3_1684_sample_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(113) is bound as output of CP function.
    -- CP-element group 114:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_4_3_1684_update_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(114) is bound as output of CP function.
    -- CP-element group 115:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: marked-predecessors 
    -- CP-element group 115: 	118 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_4_3_1684_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_4_3_1684_Sample/rr
      -- CP-element group 115: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_4_3_1684_Sample/$entry
      -- 
    rr_3509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(115), ack => RPIPE_noblock_obuf_4_3_1684_inst_req_0); -- 
    outputPort_3_Daemon_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(113) & outputPort_3_Daemon_CP_3266_elements(118);
      gj_outputPort_3_Daemon_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	117 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_4_3_1684_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_4_3_1684_Update/cr
      -- CP-element group 116: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_4_3_1684_update_start_
      -- 
    cr_3514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(116), ack => RPIPE_noblock_obuf_4_3_1684_inst_req_1); -- 
    outputPort_3_Daemon_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(117) & outputPort_3_Daemon_CP_3266_elements(114);
      gj_outputPort_3_Daemon_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	116 
    -- CP-element group 117:  members (4) 
      -- CP-element group 117: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_4_3_1684_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_4_3_1684_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_4_3_1684_Sample/ra
      -- CP-element group 117: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_4_3_1684_sample_completed__ps
      -- 
    ra_3510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_3_1684_inst_ack_0, ack => outputPort_3_Daemon_CP_3266_elements(117)); -- 
    -- CP-element group 118:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: marked-successors 
    -- CP-element group 118: 	115 
    -- CP-element group 118:  members (4) 
      -- CP-element group 118: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_4_3_1684_update_completed__ps
      -- CP-element group 118: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_4_3_1684_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_4_3_1684_Update/ca
      -- CP-element group 118: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/RPIPE_noblock_obuf_4_3_1684_update_completed_
      -- 
    ca_3515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_3_1684_inst_ack_1, ack => outputPort_3_Daemon_CP_3266_elements(118)); -- 
    -- CP-element group 119:  join  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	9 
    -- CP-element group 119: marked-predecessors 
    -- CP-element group 119: 	12 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	11 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1685_sample_start_
      -- 
    outputPort_3_Daemon_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(9) & outputPort_3_Daemon_CP_3266_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  join  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	9 
    -- CP-element group 120: marked-predecessors 
    -- CP-element group 120: 	176 
    -- CP-element group 120: 	179 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	14 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1685_update_start_
      -- 
    outputPort_3_Daemon_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(9) & outputPort_3_Daemon_CP_3266_elements(176) & outputPort_3_Daemon_CP_3266_elements(179);
      gj_outputPort_3_Daemon_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	11 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1685_sample_start__ps
      -- 
    outputPort_3_Daemon_CP_3266_elements(121) <= outputPort_3_Daemon_CP_3266_elements(11);
    -- CP-element group 122:  join  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	12 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1685_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(122) is bound as output of CP function.
    -- CP-element group 123:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	174 
    -- CP-element group 123: 	178 
    -- CP-element group 123: 	15 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1685_update_completed_
      -- CP-element group 123: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1685_update_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(123) is bound as output of CP function.
    -- CP-element group 124:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	7 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1685_loopback_trigger
      -- 
    outputPort_3_Daemon_CP_3266_elements(124) <= outputPort_3_Daemon_CP_3266_elements(7);
    -- CP-element group 125:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1685_loopback_sample_req
      -- CP-element group 125: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1685_loopback_sample_req_ps
      -- 
    phi_stmt_1685_loopback_sample_req_3526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1685_loopback_sample_req_3526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(125), ack => phi_stmt_1685_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(125) is bound as output of CP function.
    -- CP-element group 126:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	8 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1685_entry_trigger
      -- 
    outputPort_3_Daemon_CP_3266_elements(126) <= outputPort_3_Daemon_CP_3266_elements(8);
    -- CP-element group 127:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1685_entry_sample_req_ps
      -- CP-element group 127: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1685_entry_sample_req
      -- 
    phi_stmt_1685_entry_sample_req_3529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1685_entry_sample_req_3529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(127), ack => phi_stmt_1685_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(127) is bound as output of CP function.
    -- CP-element group 128:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1685_phi_mux_ack_ps
      -- CP-element group 128: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1685_phi_mux_ack
      -- 
    phi_stmt_1685_phi_mux_ack_3532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1685_ack_0, ack => outputPort_3_Daemon_CP_3266_elements(128)); -- 
    -- CP-element group 129:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (4) 
      -- CP-element group 129: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_3_1687_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_3_1687_sample_start_
      -- CP-element group 129: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_3_1687_sample_completed__ps
      -- CP-element group 129: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_3_1687_sample_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(129) is bound as output of CP function.
    -- CP-element group 130:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (2) 
      -- CP-element group 130: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_3_1687_update_start_
      -- CP-element group 130: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_3_1687_update_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(130) is bound as output of CP function.
    -- CP-element group 131:  join  transition  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	132 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_3_1687_update_completed__ps
      -- 
    outputPort_3_Daemon_CP_3266_elements(131) <= outputPort_3_Daemon_CP_3266_elements(132);
    -- CP-element group 132:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	131 
    -- CP-element group 132:  members (1) 
      -- CP-element group 132: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_3_1687_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(132) is a control-delay.
    cp_element_132_delay: control_delay_element  generic map(name => " 132_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_3266_elements(130), ack => outputPort_3_Daemon_CP_3266_elements(132), clk => clk, reset =>reset);
    -- CP-element group 133:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	135 
    -- CP-element group 133:  members (4) 
      -- CP-element group 133: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_1688_sample_start__ps
      -- CP-element group 133: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_1688_Sample/$entry
      -- CP-element group 133: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_1688_Sample/req
      -- CP-element group 133: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_1688_sample_start_
      -- 
    req_3553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(133), ack => next_active_packet_1795_1688_buf_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(133) is bound as output of CP function.
    -- CP-element group 134:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (4) 
      -- CP-element group 134: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_1688_update_start_
      -- CP-element group 134: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_1688_update_start__ps
      -- CP-element group 134: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_1688_Update/req
      -- CP-element group 134: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_1688_Update/$entry
      -- 
    req_3558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(134), ack => next_active_packet_1795_1688_buf_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(134) is bound as output of CP function.
    -- CP-element group 135:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	133 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (4) 
      -- CP-element group 135: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_1688_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_1688_sample_completed__ps
      -- CP-element group 135: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_1688_Sample/ack
      -- CP-element group 135: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_1688_Sample/$exit
      -- 
    ack_3554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_1795_1688_buf_ack_0, ack => outputPort_3_Daemon_CP_3266_elements(135)); -- 
    -- CP-element group 136:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (4) 
      -- CP-element group 136: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_1688_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_1688_update_completed__ps
      -- CP-element group 136: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_1688_Update/ack
      -- CP-element group 136: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_1688_Update/$exit
      -- 
    ack_3559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_1795_1688_buf_ack_1, ack => outputPort_3_Daemon_CP_3266_elements(136)); -- 
    -- CP-element group 137:  join  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	9 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	12 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	11 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1689_sample_start_
      -- 
    outputPort_3_Daemon_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(9) & outputPort_3_Daemon_CP_3266_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  join  transition  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	9 
    -- CP-element group 138: marked-predecessors 
    -- CP-element group 138: 	142 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	14 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1689_update_start_
      -- 
    outputPort_3_Daemon_cp_element_group_138: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_138"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(9) & outputPort_3_Daemon_CP_3266_elements(142);
      gj_outputPort_3_Daemon_cp_element_group_138 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(138), clk => clk, reset => reset); --
    end block;
    -- CP-element group 139:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	11 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1689_sample_start__ps
      -- 
    outputPort_3_Daemon_CP_3266_elements(139) <= outputPort_3_Daemon_CP_3266_elements(11);
    -- CP-element group 140:  join  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	12 
    -- CP-element group 140:  members (1) 
      -- CP-element group 140: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1689_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(140) is bound as output of CP function.
    -- CP-element group 141:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	14 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (1) 
      -- CP-element group 141: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1689_update_start__ps
      -- 
    outputPort_3_Daemon_CP_3266_elements(141) <= outputPort_3_Daemon_CP_3266_elements(14);
    -- CP-element group 142:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	15 
    -- CP-element group 142: marked-successors 
    -- CP-element group 142: 	138 
    -- CP-element group 142:  members (2) 
      -- CP-element group 142: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1689_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1689_update_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(142) is bound as output of CP function.
    -- CP-element group 143:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	7 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1689_loopback_trigger
      -- 
    outputPort_3_Daemon_CP_3266_elements(143) <= outputPort_3_Daemon_CP_3266_elements(7);
    -- CP-element group 144:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (2) 
      -- CP-element group 144: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1689_loopback_sample_req
      -- CP-element group 144: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1689_loopback_sample_req_ps
      -- 
    phi_stmt_1689_loopback_sample_req_3570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1689_loopback_sample_req_3570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(144), ack => phi_stmt_1689_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(144) is bound as output of CP function.
    -- CP-element group 145:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	8 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (1) 
      -- CP-element group 145: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1689_entry_trigger
      -- 
    outputPort_3_Daemon_CP_3266_elements(145) <= outputPort_3_Daemon_CP_3266_elements(8);
    -- CP-element group 146:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (2) 
      -- CP-element group 146: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1689_entry_sample_req
      -- CP-element group 146: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1689_entry_sample_req_ps
      -- 
    phi_stmt_1689_entry_sample_req_3573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1689_entry_sample_req_3573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(146), ack => phi_stmt_1689_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(146) is bound as output of CP function.
    -- CP-element group 147:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (2) 
      -- CP-element group 147: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1689_phi_mux_ack
      -- CP-element group 147: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1689_phi_mux_ack_ps
      -- 
    phi_stmt_1689_phi_mux_ack_3576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1689_ack_0, ack => outputPort_3_Daemon_CP_3266_elements(147)); -- 
    -- CP-element group 148:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (4) 
      -- CP-element group 148: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_8_1691_sample_start__ps
      -- CP-element group 148: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_8_1691_sample_completed__ps
      -- CP-element group 148: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_8_1691_sample_start_
      -- CP-element group 148: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_8_1691_sample_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(148) is bound as output of CP function.
    -- CP-element group 149:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	151 
    -- CP-element group 149:  members (2) 
      -- CP-element group 149: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_8_1691_update_start__ps
      -- CP-element group 149: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_8_1691_update_start_
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(149) is bound as output of CP function.
    -- CP-element group 150:  join  transition  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	151 
    -- CP-element group 150: successors 
    -- CP-element group 150:  members (1) 
      -- CP-element group 150: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_8_1691_update_completed__ps
      -- 
    outputPort_3_Daemon_CP_3266_elements(150) <= outputPort_3_Daemon_CP_3266_elements(151);
    -- CP-element group 151:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	149 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	150 
    -- CP-element group 151:  members (1) 
      -- CP-element group 151: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_8_1691_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(151) is a control-delay.
    cp_element_151_delay: control_delay_element  generic map(name => " 151_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_3266_elements(149), ack => outputPort_3_Daemon_CP_3266_elements(151), clk => clk, reset =>reset);
    -- CP-element group 152:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (4) 
      -- CP-element group 152: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_length_1692_sample_start__ps
      -- CP-element group 152: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_length_1692_sample_start_
      -- CP-element group 152: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_length_1692_Sample/$entry
      -- CP-element group 152: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_length_1692_Sample/req
      -- 
    req_3597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(152), ack => next_active_packet_length_1840_1692_buf_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(152) is bound as output of CP function.
    -- CP-element group 153:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	155 
    -- CP-element group 153:  members (4) 
      -- CP-element group 153: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_length_1692_update_start__ps
      -- CP-element group 153: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_length_1692_update_start_
      -- CP-element group 153: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_length_1692_Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_length_1692_Update/req
      -- 
    req_3602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(153), ack => next_active_packet_length_1840_1692_buf_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(153) is bound as output of CP function.
    -- CP-element group 154:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	152 
    -- CP-element group 154: successors 
    -- CP-element group 154:  members (4) 
      -- CP-element group 154: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_length_1692_sample_completed__ps
      -- CP-element group 154: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_length_1692_sample_completed_
      -- CP-element group 154: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_length_1692_Sample/$exit
      -- CP-element group 154: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_length_1692_Sample/ack
      -- 
    ack_3598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_length_1840_1692_buf_ack_0, ack => outputPort_3_Daemon_CP_3266_elements(154)); -- 
    -- CP-element group 155:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	153 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (4) 
      -- CP-element group 155: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_length_1692_update_completed__ps
      -- CP-element group 155: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_length_1692_update_completed_
      -- CP-element group 155: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_length_1692_Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_active_packet_length_1692_Update/ack
      -- 
    ack_3603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_length_1840_1692_buf_ack_1, ack => outputPort_3_Daemon_CP_3266_elements(155)); -- 
    -- CP-element group 156:  join  transition  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	9 
    -- CP-element group 156: marked-predecessors 
    -- CP-element group 156: 	12 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	11 
    -- CP-element group 156:  members (1) 
      -- CP-element group 156: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1693_sample_start_
      -- 
    outputPort_3_Daemon_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(9) & outputPort_3_Daemon_CP_3266_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  join  transition  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	9 
    -- CP-element group 157: marked-predecessors 
    -- CP-element group 157: 	176 
    -- CP-element group 157: 	179 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	14 
    -- CP-element group 157:  members (1) 
      -- CP-element group 157: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1693_update_start_
      -- 
    outputPort_3_Daemon_cp_element_group_157: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_157"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(9) & outputPort_3_Daemon_CP_3266_elements(176) & outputPort_3_Daemon_CP_3266_elements(179);
      gj_outputPort_3_Daemon_cp_element_group_157 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(157), clk => clk, reset => reset); --
    end block;
    -- CP-element group 158:  join  transition  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	12 
    -- CP-element group 158:  members (1) 
      -- CP-element group 158: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1693_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(158) is bound as output of CP function.
    -- CP-element group 159:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	14 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (1) 
      -- CP-element group 159: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1693_update_start__ps
      -- 
    outputPort_3_Daemon_CP_3266_elements(159) <= outputPort_3_Daemon_CP_3266_elements(14);
    -- CP-element group 160:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	174 
    -- CP-element group 160: 	178 
    -- CP-element group 160: 	15 
    -- CP-element group 160:  members (2) 
      -- CP-element group 160: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1693_update_completed_
      -- CP-element group 160: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1693_update_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(160) is bound as output of CP function.
    -- CP-element group 161:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	7 
    -- CP-element group 161: successors 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1693_loopback_trigger
      -- 
    outputPort_3_Daemon_CP_3266_elements(161) <= outputPort_3_Daemon_CP_3266_elements(7);
    -- CP-element group 162:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (2) 
      -- CP-element group 162: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1693_loopback_sample_req
      -- CP-element group 162: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1693_loopback_sample_req_ps
      -- 
    phi_stmt_1693_loopback_sample_req_3614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1693_loopback_sample_req_3614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(162), ack => phi_stmt_1693_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(162) is bound as output of CP function.
    -- CP-element group 163:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	8 
    -- CP-element group 163: successors 
    -- CP-element group 163:  members (1) 
      -- CP-element group 163: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1693_entry_trigger
      -- 
    outputPort_3_Daemon_CP_3266_elements(163) <= outputPort_3_Daemon_CP_3266_elements(8);
    -- CP-element group 164:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (2) 
      -- CP-element group 164: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1693_entry_sample_req
      -- CP-element group 164: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1693_entry_sample_req_ps
      -- 
    phi_stmt_1693_entry_sample_req_3617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1693_entry_sample_req_3617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(164), ack => phi_stmt_1693_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(164) is bound as output of CP function.
    -- CP-element group 165:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: successors 
    -- CP-element group 165:  members (2) 
      -- CP-element group 165: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1693_phi_mux_ack
      -- CP-element group 165: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/phi_stmt_1693_phi_mux_ack_ps
      -- 
    phi_stmt_1693_phi_mux_ack_3620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1693_ack_0, ack => outputPort_3_Daemon_CP_3266_elements(165)); -- 
    -- CP-element group 166:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	168 
    -- CP-element group 166:  members (4) 
      -- CP-element group 166: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_priority_index_1695_sample_start__ps
      -- CP-element group 166: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_priority_index_1695_sample_start_
      -- CP-element group 166: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_priority_index_1695_Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_priority_index_1695_Sample/req
      -- 
    req_3633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(166), ack => next_priority_index_1795_1695_buf_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(166) is bound as output of CP function.
    -- CP-element group 167:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (4) 
      -- CP-element group 167: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_priority_index_1695_update_start__ps
      -- CP-element group 167: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_priority_index_1695_update_start_
      -- CP-element group 167: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_priority_index_1695_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_priority_index_1695_Update/req
      -- 
    req_3638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(167), ack => next_priority_index_1795_1695_buf_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(167) is bound as output of CP function.
    -- CP-element group 168:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	166 
    -- CP-element group 168: successors 
    -- CP-element group 168:  members (4) 
      -- CP-element group 168: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_priority_index_1695_sample_completed__ps
      -- CP-element group 168: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_priority_index_1695_sample_completed_
      -- CP-element group 168: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_priority_index_1695_Sample/$exit
      -- CP-element group 168: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_priority_index_1695_Sample/ack
      -- 
    ack_3634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_priority_index_1795_1695_buf_ack_0, ack => outputPort_3_Daemon_CP_3266_elements(168)); -- 
    -- CP-element group 169:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169:  members (4) 
      -- CP-element group 169: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_priority_index_1695_update_completed__ps
      -- CP-element group 169: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_priority_index_1695_update_completed_
      -- CP-element group 169: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_priority_index_1695_Update/$exit
      -- CP-element group 169: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_next_priority_index_1695_Update/ack
      -- 
    ack_3639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_priority_index_1795_1695_buf_ack_1, ack => outputPort_3_Daemon_CP_3266_elements(169)); -- 
    -- CP-element group 170:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: successors 
    -- CP-element group 170:  members (4) 
      -- CP-element group 170: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_2_1696_sample_start__ps
      -- CP-element group 170: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_2_1696_sample_completed__ps
      -- CP-element group 170: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_2_1696_sample_start_
      -- CP-element group 170: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_2_1696_sample_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(170) is bound as output of CP function.
    -- CP-element group 171:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (2) 
      -- CP-element group 171: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_2_1696_update_start__ps
      -- CP-element group 171: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_2_1696_update_start_
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(171) is bound as output of CP function.
    -- CP-element group 172:  join  transition  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	173 
    -- CP-element group 172: successors 
    -- CP-element group 172:  members (1) 
      -- CP-element group 172: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_2_1696_update_completed__ps
      -- 
    outputPort_3_Daemon_CP_3266_elements(172) <= outputPort_3_Daemon_CP_3266_elements(173);
    -- CP-element group 173:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	172 
    -- CP-element group 173:  members (1) 
      -- CP-element group 173: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/R_ZERO_2_1696_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(173) is a control-delay.
    cp_element_173_delay: control_delay_element  generic map(name => " 173_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_3266_elements(171), ack => outputPort_3_Daemon_CP_3266_elements(173), clk => clk, reset =>reset);
    -- CP-element group 174:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	123 
    -- CP-element group 174: 	160 
    -- CP-element group 174: 	82 
    -- CP-element group 174: 	103 
    -- CP-element group 174: 	21 
    -- CP-element group 174: 	40 
    -- CP-element group 174: 	61 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	176 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/call_stmt_1724_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/call_stmt_1724_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/call_stmt_1724_Sample/crr
      -- 
    crr_3656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(174), ack => call_stmt_1724_call_req_0); -- 
    outputPort_3_Daemon_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(123) & outputPort_3_Daemon_CP_3266_elements(160) & outputPort_3_Daemon_CP_3266_elements(82) & outputPort_3_Daemon_CP_3266_elements(103) & outputPort_3_Daemon_CP_3266_elements(21) & outputPort_3_Daemon_CP_3266_elements(40) & outputPort_3_Daemon_CP_3266_elements(61);
      gj_outputPort_3_Daemon_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: marked-predecessors 
    -- CP-element group 175: 	177 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	177 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/call_stmt_1724_update_start_
      -- CP-element group 175: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/call_stmt_1724_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/call_stmt_1724_Update/ccr
      -- 
    ccr_3661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(175), ack => call_stmt_1724_call_req_1); -- 
    outputPort_3_Daemon_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= outputPort_3_Daemon_CP_3266_elements(177);
      gj_outputPort_3_Daemon_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	174 
    -- CP-element group 176: successors 
    -- CP-element group 176: marked-successors 
    -- CP-element group 176: 	157 
    -- CP-element group 176: 	120 
    -- CP-element group 176: 	78 
    -- CP-element group 176: 	99 
    -- CP-element group 176: 	17 
    -- CP-element group 176: 	36 
    -- CP-element group 176: 	57 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/call_stmt_1724_sample_completed_
      -- CP-element group 176: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/call_stmt_1724_Sample/$exit
      -- CP-element group 176: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/call_stmt_1724_Sample/cra
      -- 
    cra_3657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1724_call_ack_0, ack => outputPort_3_Daemon_CP_3266_elements(176)); -- 
    -- CP-element group 177:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	182 
    -- CP-element group 177: marked-successors 
    -- CP-element group 177: 	175 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/call_stmt_1724_update_completed_
      -- CP-element group 177: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/call_stmt_1724_Update/$exit
      -- CP-element group 177: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/call_stmt_1724_Update/cca
      -- 
    cca_3662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1724_call_ack_1, ack => outputPort_3_Daemon_CP_3266_elements(177)); -- 
    -- CP-element group 178:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	123 
    -- CP-element group 178: 	160 
    -- CP-element group 178: 	82 
    -- CP-element group 178: 	103 
    -- CP-element group 178: 	21 
    -- CP-element group 178: 	40 
    -- CP-element group 178: 	61 
    -- CP-element group 178: marked-predecessors 
    -- CP-element group 178: 	180 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/WPIPE_out_data_3_1949_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/WPIPE_out_data_3_1949_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/WPIPE_out_data_3_1949_Sample/req
      -- 
    req_3670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(178), ack => WPIPE_out_data_3_1949_inst_req_0); -- 
    outputPort_3_Daemon_cp_element_group_178: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_178"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(123) & outputPort_3_Daemon_CP_3266_elements(160) & outputPort_3_Daemon_CP_3266_elements(82) & outputPort_3_Daemon_CP_3266_elements(103) & outputPort_3_Daemon_CP_3266_elements(21) & outputPort_3_Daemon_CP_3266_elements(40) & outputPort_3_Daemon_CP_3266_elements(61) & outputPort_3_Daemon_CP_3266_elements(180);
      gj_outputPort_3_Daemon_cp_element_group_178 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(178), clk => clk, reset => reset); --
    end block;
    -- CP-element group 179:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179: marked-successors 
    -- CP-element group 179: 	157 
    -- CP-element group 179: 	120 
    -- CP-element group 179: 	78 
    -- CP-element group 179: 	99 
    -- CP-element group 179: 	17 
    -- CP-element group 179: 	36 
    -- CP-element group 179: 	57 
    -- CP-element group 179:  members (6) 
      -- CP-element group 179: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/WPIPE_out_data_3_1949_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/WPIPE_out_data_3_1949_update_start_
      -- CP-element group 179: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/WPIPE_out_data_3_1949_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/WPIPE_out_data_3_1949_Sample/ack
      -- CP-element group 179: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/WPIPE_out_data_3_1949_Update/$entry
      -- CP-element group 179: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/WPIPE_out_data_3_1949_Update/req
      -- 
    ack_3671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_3_1949_inst_ack_0, ack => outputPort_3_Daemon_CP_3266_elements(179)); -- 
    req_3675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_3266_elements(179), ack => WPIPE_out_data_3_1949_inst_req_1); -- 
    -- CP-element group 180:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	182 
    -- CP-element group 180: marked-successors 
    -- CP-element group 180: 	178 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/WPIPE_out_data_3_1949_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/WPIPE_out_data_3_1949_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/WPIPE_out_data_3_1949_Update/ack
      -- 
    ack_3676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_3_1949_inst_ack_1, ack => outputPort_3_Daemon_CP_3266_elements(180)); -- 
    -- CP-element group 181:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	9 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	10 
    -- CP-element group 181:  members (1) 
      -- CP-element group 181: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group outputPort_3_Daemon_CP_3266_elements(181) is a control-delay.
    cp_element_181_delay: control_delay_element  generic map(name => " 181_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_3266_elements(9), ack => outputPort_3_Daemon_CP_3266_elements(181), clk => clk, reset =>reset);
    -- CP-element group 182:  join  transition  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	177 
    -- CP-element group 182: 	180 
    -- CP-element group 182: 	12 
    -- CP-element group 182: 	13 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	6 
    -- CP-element group 182:  members (1) 
      -- CP-element group 182: 	 branch_block_stmt_1658/do_while_stmt_1659/do_while_stmt_1659_loop_body/$exit
      -- 
    outputPort_3_Daemon_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 7,2 => 7,3 => 7);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_3266_elements(177) & outputPort_3_Daemon_CP_3266_elements(180) & outputPort_3_Daemon_CP_3266_elements(12) & outputPort_3_Daemon_CP_3266_elements(13);
      gj_outputPort_3_Daemon_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  transition  input  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	5 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (2) 
      -- CP-element group 183: 	 branch_block_stmt_1658/do_while_stmt_1659/loop_exit/$exit
      -- CP-element group 183: 	 branch_block_stmt_1658/do_while_stmt_1659/loop_exit/ack
      -- 
    ack_3681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1659_branch_ack_0, ack => outputPort_3_Daemon_CP_3266_elements(183)); -- 
    -- CP-element group 184:  transition  input  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	5 
    -- CP-element group 184: successors 
    -- CP-element group 184:  members (2) 
      -- CP-element group 184: 	 branch_block_stmt_1658/do_while_stmt_1659/loop_taken/$exit
      -- CP-element group 184: 	 branch_block_stmt_1658/do_while_stmt_1659/loop_taken/ack
      -- 
    ack_3685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1659_branch_ack_1, ack => outputPort_3_Daemon_CP_3266_elements(184)); -- 
    -- CP-element group 185:  transition  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	3 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	1 
    -- CP-element group 185:  members (1) 
      -- CP-element group 185: 	 branch_block_stmt_1658/do_while_stmt_1659/$exit
      -- 
    outputPort_3_Daemon_CP_3266_elements(185) <= outputPort_3_Daemon_CP_3266_elements(3);
    outputPort_3_Daemon_do_while_stmt_1659_terminator_3686: loop_terminator -- 
      generic map (name => " outputPort_3_Daemon_do_while_stmt_1659_terminator_3686", max_iterations_in_flight =>7) 
      port map(loop_body_exit => outputPort_3_Daemon_CP_3266_elements(6),loop_continue => outputPort_3_Daemon_CP_3266_elements(184),loop_terminate => outputPort_3_Daemon_CP_3266_elements(183),loop_back => outputPort_3_Daemon_CP_3266_elements(4),loop_exit => outputPort_3_Daemon_CP_3266_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1661_phi_seq_3340_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_3_Daemon_CP_3266_elements(24);
      outputPort_3_Daemon_CP_3266_elements(27)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_3_Daemon_CP_3266_elements(27);
      outputPort_3_Daemon_CP_3266_elements(28)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_3_Daemon_CP_3266_elements(29);
      outputPort_3_Daemon_CP_3266_elements(25) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_3_Daemon_CP_3266_elements(22);
      outputPort_3_Daemon_CP_3266_elements(31)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_3_Daemon_CP_3266_elements(33);
      outputPort_3_Daemon_CP_3266_elements(32)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_3_Daemon_CP_3266_elements(34);
      outputPort_3_Daemon_CP_3266_elements(23) <= phi_mux_reqs(1);
      phi_stmt_1661_phi_seq_3340 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1661_phi_seq_3340") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_3_Daemon_CP_3266_elements(18), 
          phi_sample_ack => outputPort_3_Daemon_CP_3266_elements(19), 
          phi_update_req => outputPort_3_Daemon_CP_3266_elements(20), 
          phi_update_ack => outputPort_3_Daemon_CP_3266_elements(21), 
          phi_mux_ack => outputPort_3_Daemon_CP_3266_elements(26), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1665_phi_seq_3384_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_3_Daemon_CP_3266_elements(43);
      outputPort_3_Daemon_CP_3266_elements(46)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_3_Daemon_CP_3266_elements(46);
      outputPort_3_Daemon_CP_3266_elements(47)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_3_Daemon_CP_3266_elements(48);
      outputPort_3_Daemon_CP_3266_elements(44) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_3_Daemon_CP_3266_elements(41);
      outputPort_3_Daemon_CP_3266_elements(50)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_3_Daemon_CP_3266_elements(54);
      outputPort_3_Daemon_CP_3266_elements(51)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_3_Daemon_CP_3266_elements(55);
      outputPort_3_Daemon_CP_3266_elements(42) <= phi_mux_reqs(1);
      phi_stmt_1665_phi_seq_3384 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1665_phi_seq_3384") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_3_Daemon_CP_3266_elements(37), 
          phi_sample_ack => outputPort_3_Daemon_CP_3266_elements(38), 
          phi_update_req => outputPort_3_Daemon_CP_3266_elements(39), 
          phi_update_ack => outputPort_3_Daemon_CP_3266_elements(40), 
          phi_mux_ack => outputPort_3_Daemon_CP_3266_elements(45), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1670_phi_seq_3428_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_3_Daemon_CP_3266_elements(64);
      outputPort_3_Daemon_CP_3266_elements(67)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_3_Daemon_CP_3266_elements(67);
      outputPort_3_Daemon_CP_3266_elements(68)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_3_Daemon_CP_3266_elements(69);
      outputPort_3_Daemon_CP_3266_elements(65) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_3_Daemon_CP_3266_elements(62);
      outputPort_3_Daemon_CP_3266_elements(71)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_3_Daemon_CP_3266_elements(75);
      outputPort_3_Daemon_CP_3266_elements(72)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_3_Daemon_CP_3266_elements(76);
      outputPort_3_Daemon_CP_3266_elements(63) <= phi_mux_reqs(1);
      phi_stmt_1670_phi_seq_3428 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1670_phi_seq_3428") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_3_Daemon_CP_3266_elements(58), 
          phi_sample_ack => outputPort_3_Daemon_CP_3266_elements(59), 
          phi_update_req => outputPort_3_Daemon_CP_3266_elements(60), 
          phi_update_ack => outputPort_3_Daemon_CP_3266_elements(61), 
          phi_mux_ack => outputPort_3_Daemon_CP_3266_elements(66), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1675_phi_seq_3472_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_3_Daemon_CP_3266_elements(85);
      outputPort_3_Daemon_CP_3266_elements(88)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_3_Daemon_CP_3266_elements(88);
      outputPort_3_Daemon_CP_3266_elements(89)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_3_Daemon_CP_3266_elements(90);
      outputPort_3_Daemon_CP_3266_elements(86) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_3_Daemon_CP_3266_elements(83);
      outputPort_3_Daemon_CP_3266_elements(92)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_3_Daemon_CP_3266_elements(96);
      outputPort_3_Daemon_CP_3266_elements(93)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_3_Daemon_CP_3266_elements(97);
      outputPort_3_Daemon_CP_3266_elements(84) <= phi_mux_reqs(1);
      phi_stmt_1675_phi_seq_3472 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1675_phi_seq_3472") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_3_Daemon_CP_3266_elements(79), 
          phi_sample_ack => outputPort_3_Daemon_CP_3266_elements(80), 
          phi_update_req => outputPort_3_Daemon_CP_3266_elements(81), 
          phi_update_ack => outputPort_3_Daemon_CP_3266_elements(82), 
          phi_mux_ack => outputPort_3_Daemon_CP_3266_elements(87), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1680_phi_seq_3516_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_3_Daemon_CP_3266_elements(106);
      outputPort_3_Daemon_CP_3266_elements(109)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_3_Daemon_CP_3266_elements(109);
      outputPort_3_Daemon_CP_3266_elements(110)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_3_Daemon_CP_3266_elements(111);
      outputPort_3_Daemon_CP_3266_elements(107) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_3_Daemon_CP_3266_elements(104);
      outputPort_3_Daemon_CP_3266_elements(113)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_3_Daemon_CP_3266_elements(117);
      outputPort_3_Daemon_CP_3266_elements(114)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_3_Daemon_CP_3266_elements(118);
      outputPort_3_Daemon_CP_3266_elements(105) <= phi_mux_reqs(1);
      phi_stmt_1680_phi_seq_3516 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1680_phi_seq_3516") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_3_Daemon_CP_3266_elements(100), 
          phi_sample_ack => outputPort_3_Daemon_CP_3266_elements(101), 
          phi_update_req => outputPort_3_Daemon_CP_3266_elements(102), 
          phi_update_ack => outputPort_3_Daemon_CP_3266_elements(103), 
          phi_mux_ack => outputPort_3_Daemon_CP_3266_elements(108), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1685_phi_seq_3560_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_3_Daemon_CP_3266_elements(126);
      outputPort_3_Daemon_CP_3266_elements(129)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_3_Daemon_CP_3266_elements(129);
      outputPort_3_Daemon_CP_3266_elements(130)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_3_Daemon_CP_3266_elements(131);
      outputPort_3_Daemon_CP_3266_elements(127) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_3_Daemon_CP_3266_elements(124);
      outputPort_3_Daemon_CP_3266_elements(133)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_3_Daemon_CP_3266_elements(135);
      outputPort_3_Daemon_CP_3266_elements(134)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_3_Daemon_CP_3266_elements(136);
      outputPort_3_Daemon_CP_3266_elements(125) <= phi_mux_reqs(1);
      phi_stmt_1685_phi_seq_3560 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1685_phi_seq_3560") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_3_Daemon_CP_3266_elements(121), 
          phi_sample_ack => outputPort_3_Daemon_CP_3266_elements(122), 
          phi_update_req => outputPort_3_Daemon_CP_3266_elements(14), 
          phi_update_ack => outputPort_3_Daemon_CP_3266_elements(123), 
          phi_mux_ack => outputPort_3_Daemon_CP_3266_elements(128), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1689_phi_seq_3604_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_3_Daemon_CP_3266_elements(145);
      outputPort_3_Daemon_CP_3266_elements(148)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_3_Daemon_CP_3266_elements(148);
      outputPort_3_Daemon_CP_3266_elements(149)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_3_Daemon_CP_3266_elements(150);
      outputPort_3_Daemon_CP_3266_elements(146) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_3_Daemon_CP_3266_elements(143);
      outputPort_3_Daemon_CP_3266_elements(152)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_3_Daemon_CP_3266_elements(154);
      outputPort_3_Daemon_CP_3266_elements(153)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_3_Daemon_CP_3266_elements(155);
      outputPort_3_Daemon_CP_3266_elements(144) <= phi_mux_reqs(1);
      phi_stmt_1689_phi_seq_3604 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1689_phi_seq_3604") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_3_Daemon_CP_3266_elements(139), 
          phi_sample_ack => outputPort_3_Daemon_CP_3266_elements(140), 
          phi_update_req => outputPort_3_Daemon_CP_3266_elements(141), 
          phi_update_ack => outputPort_3_Daemon_CP_3266_elements(142), 
          phi_mux_ack => outputPort_3_Daemon_CP_3266_elements(147), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1693_phi_seq_3648_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_3_Daemon_CP_3266_elements(161);
      outputPort_3_Daemon_CP_3266_elements(166)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_3_Daemon_CP_3266_elements(168);
      outputPort_3_Daemon_CP_3266_elements(167)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_3_Daemon_CP_3266_elements(169);
      outputPort_3_Daemon_CP_3266_elements(162) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_3_Daemon_CP_3266_elements(163);
      outputPort_3_Daemon_CP_3266_elements(170)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_3_Daemon_CP_3266_elements(170);
      outputPort_3_Daemon_CP_3266_elements(171)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_3_Daemon_CP_3266_elements(172);
      outputPort_3_Daemon_CP_3266_elements(164) <= phi_mux_reqs(1);
      phi_stmt_1693_phi_seq_3648 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1693_phi_seq_3648") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_3_Daemon_CP_3266_elements(11), 
          phi_sample_ack => outputPort_3_Daemon_CP_3266_elements(158), 
          phi_update_req => outputPort_3_Daemon_CP_3266_elements(159), 
          phi_update_ack => outputPort_3_Daemon_CP_3266_elements(160), 
          phi_mux_ack => outputPort_3_Daemon_CP_3266_elements(165), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3291_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= outputPort_3_Daemon_CP_3266_elements(7);
        preds(1)  <= outputPort_3_Daemon_CP_3266_elements(8);
        entry_tmerge_3291 : transition_merge -- 
          generic map(name => " entry_tmerge_3291")
          port map (preds => preds, symbol_out => outputPort_3_Daemon_CP_3266_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal EQ_u3_u1_1760_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1766_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1773_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1779_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1809_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1816_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1824_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1831_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1859_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1867_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1875_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1883_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1889_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1896_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1904_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1911_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1922_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1928_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1935_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1941_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_1802_wire : std_logic_vector(0 downto 0);
    signal MUX_1702_wire : std_logic_vector(7 downto 0);
    signal MUX_1706_wire : std_logic_vector(7 downto 0);
    signal MUX_1711_wire : std_logic_vector(7 downto 0);
    signal MUX_1715_wire : std_logic_vector(7 downto 0);
    signal MUX_1763_wire : std_logic_vector(0 downto 0);
    signal MUX_1769_wire : std_logic_vector(0 downto 0);
    signal MUX_1776_wire : std_logic_vector(0 downto 0);
    signal MUX_1782_wire : std_logic_vector(0 downto 0);
    signal MUX_1813_wire : std_logic_vector(7 downto 0);
    signal MUX_1820_wire : std_logic_vector(7 downto 0);
    signal MUX_1828_wire : std_logic_vector(7 downto 0);
    signal MUX_1835_wire : std_logic_vector(7 downto 0);
    signal MUX_1851_wire : std_logic_vector(7 downto 0);
    signal MUX_1893_wire : std_logic_vector(31 downto 0);
    signal MUX_1900_wire : std_logic_vector(31 downto 0);
    signal MUX_1908_wire : std_logic_vector(31 downto 0);
    signal MUX_1915_wire : std_logic_vector(31 downto 0);
    signal MUX_1925_wire : std_logic_vector(0 downto 0);
    signal MUX_1931_wire : std_logic_vector(0 downto 0);
    signal MUX_1938_wire : std_logic_vector(0 downto 0);
    signal MUX_1944_wire : std_logic_vector(0 downto 0);
    signal NEQ_u3_u1_1799_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1856_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1864_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1872_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1880_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1770_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1783_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1932_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1945_wire : std_logic_vector(0 downto 0);
    signal OR_u32_u32_1901_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_1916_wire : std_logic_vector(31 downto 0);
    signal OR_u8_u8_1707_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_1716_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_1821_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_1836_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_1837_wire : std_logic_vector(7 downto 0);
    signal RPIPE_noblock_obuf_1_3_1669_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_2_3_1674_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_3_3_1679_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_4_3_1684_wire : std_logic_vector(32 downto 0);
    signal R_ZERO_2_1696_wire_constant : std_logic_vector(1 downto 0);
    signal R_ZERO_33_1667_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1672_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1677_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1682_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_3_1687_wire_constant : std_logic_vector(2 downto 0);
    signal R_ZERO_8_1663_wire_constant : std_logic_vector(7 downto 0);
    signal R_ZERO_8_1691_wire_constant : std_logic_vector(7 downto 0);
    signal SUB_u8_u8_1845_wire : std_logic_vector(7 downto 0);
    signal SUB_u8_u8_1849_wire : std_logic_vector(7 downto 0);
    signal active_packet_1685 : std_logic_vector(2 downto 0);
    signal active_packet_length_1689 : std_logic_vector(7 downto 0);
    signal continue_1724 : std_logic_vector(0 downto 0);
    signal data_to_out_1918 : std_logic_vector(31 downto 0);
    signal down_counter_1661 : std_logic_vector(7 downto 0);
    signal konst_1700_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1701_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1704_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1705_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1709_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1710_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1713_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1714_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1720_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1727_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1732_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1737_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1742_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1759_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1762_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1765_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1768_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1772_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1775_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1778_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1781_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1798_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1801_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1808_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1812_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1815_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1819_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1823_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1827_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1830_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1834_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1844_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1848_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1858_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1866_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1874_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1882_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1888_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1892_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1895_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1899_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1903_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1907_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1910_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1914_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1921_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1924_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1927_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1930_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1934_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1937_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1940_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1943_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1962_wire_constant : std_logic_vector(0 downto 0);
    signal next_active_packet_1795 : std_logic_vector(2 downto 0);
    signal next_active_packet_1795_1688_buffered : std_logic_vector(2 downto 0);
    signal next_active_packet_length_1840 : std_logic_vector(7 downto 0);
    signal next_active_packet_length_1840_1692_buffered : std_logic_vector(7 downto 0);
    signal next_down_counter_1853 : std_logic_vector(7 downto 0);
    signal next_down_counter_1853_1664_buffered : std_logic_vector(7 downto 0);
    signal next_priority_index_1795 : std_logic_vector(1 downto 0);
    signal next_priority_index_1795_1695_buffered : std_logic_vector(1 downto 0);
    signal p1_valid_1729 : std_logic_vector(0 downto 0);
    signal p2_valid_1734 : std_logic_vector(0 downto 0);
    signal p3_valid_1739 : std_logic_vector(0 downto 0);
    signal p4_valid_1744 : std_logic_vector(0 downto 0);
    signal pkt_1_e_word_1665 : std_logic_vector(32 downto 0);
    signal pkt_2_e_word_1670 : std_logic_vector(32 downto 0);
    signal pkt_3_e_word_1675 : std_logic_vector(32 downto 0);
    signal pkt_4_e_word_1680 : std_logic_vector(32 downto 0);
    signal priority_index_1693 : std_logic_vector(1 downto 0);
    signal read_from_1_1861 : std_logic_vector(0 downto 0);
    signal read_from_2_1869 : std_logic_vector(0 downto 0);
    signal read_from_3_1877 : std_logic_vector(0 downto 0);
    signal read_from_4_1885 : std_logic_vector(0 downto 0);
    signal send_flag_1947 : std_logic_vector(0 downto 0);
    signal senderPort_1718 : std_logic_vector(7 downto 0);
    signal slice_1811_wire : std_logic_vector(7 downto 0);
    signal slice_1818_wire : std_logic_vector(7 downto 0);
    signal slice_1826_wire : std_logic_vector(7 downto 0);
    signal slice_1833_wire : std_logic_vector(7 downto 0);
    signal slice_1891_wire : std_logic_vector(31 downto 0);
    signal slice_1898_wire : std_logic_vector(31 downto 0);
    signal slice_1906_wire : std_logic_vector(31 downto 0);
    signal slice_1913_wire : std_logic_vector(31 downto 0);
    signal started_new_packet_1804 : std_logic_vector(0 downto 0);
    signal type_cast_1722_wire_constant : std_logic_vector(0 downto 0);
    signal valid_active_pkt_word_read_1785 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_ZERO_2_1696_wire_constant <= "00";
    R_ZERO_33_1667_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1672_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1677_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1682_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_3_1687_wire_constant <= "000";
    R_ZERO_8_1663_wire_constant <= "00000000";
    R_ZERO_8_1691_wire_constant <= "00000000";
    konst_1700_wire_constant <= "00000000";
    konst_1701_wire_constant <= "00000000";
    konst_1704_wire_constant <= "00000001";
    konst_1705_wire_constant <= "00000000";
    konst_1709_wire_constant <= "00000010";
    konst_1710_wire_constant <= "00000000";
    konst_1713_wire_constant <= "00000011";
    konst_1714_wire_constant <= "00000000";
    konst_1720_wire_constant <= "00000010";
    konst_1727_wire_constant <= "000000000000000000000000000100000";
    konst_1732_wire_constant <= "000000000000000000000000000100000";
    konst_1737_wire_constant <= "000000000000000000000000000100000";
    konst_1742_wire_constant <= "000000000000000000000000000100000";
    konst_1759_wire_constant <= "001";
    konst_1762_wire_constant <= "0";
    konst_1765_wire_constant <= "010";
    konst_1768_wire_constant <= "0";
    konst_1772_wire_constant <= "011";
    konst_1775_wire_constant <= "0";
    konst_1778_wire_constant <= "100";
    konst_1781_wire_constant <= "0";
    konst_1798_wire_constant <= "000";
    konst_1801_wire_constant <= "00000000";
    konst_1808_wire_constant <= "001";
    konst_1812_wire_constant <= "00000000";
    konst_1815_wire_constant <= "010";
    konst_1819_wire_constant <= "00000000";
    konst_1823_wire_constant <= "011";
    konst_1827_wire_constant <= "00000000";
    konst_1830_wire_constant <= "100";
    konst_1834_wire_constant <= "00000000";
    konst_1844_wire_constant <= "00000001";
    konst_1848_wire_constant <= "00000001";
    konst_1858_wire_constant <= "001";
    konst_1866_wire_constant <= "010";
    konst_1874_wire_constant <= "011";
    konst_1882_wire_constant <= "100";
    konst_1888_wire_constant <= "001";
    konst_1892_wire_constant <= "00000000000000000000000000000000";
    konst_1895_wire_constant <= "010";
    konst_1899_wire_constant <= "00000000000000000000000000000000";
    konst_1903_wire_constant <= "011";
    konst_1907_wire_constant <= "00000000000000000000000000000000";
    konst_1910_wire_constant <= "100";
    konst_1914_wire_constant <= "00000000000000000000000000000000";
    konst_1921_wire_constant <= "001";
    konst_1924_wire_constant <= "0";
    konst_1927_wire_constant <= "010";
    konst_1930_wire_constant <= "0";
    konst_1934_wire_constant <= "011";
    konst_1937_wire_constant <= "0";
    konst_1940_wire_constant <= "100";
    konst_1943_wire_constant <= "0";
    konst_1962_wire_constant <= "1";
    type_cast_1722_wire_constant <= "0";
    phi_stmt_1661: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_8_1663_wire_constant & next_down_counter_1853_1664_buffered;
      req <= phi_stmt_1661_req_0 & phi_stmt_1661_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1661",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1661_ack_0,
          idata => idata,
          odata => down_counter_1661,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1661
    phi_stmt_1665: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1667_wire_constant & RPIPE_noblock_obuf_1_3_1669_wire;
      req <= phi_stmt_1665_req_0 & phi_stmt_1665_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1665",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1665_ack_0,
          idata => idata,
          odata => pkt_1_e_word_1665,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1665
    phi_stmt_1670: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1672_wire_constant & RPIPE_noblock_obuf_2_3_1674_wire;
      req <= phi_stmt_1670_req_0 & phi_stmt_1670_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1670",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1670_ack_0,
          idata => idata,
          odata => pkt_2_e_word_1670,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1670
    phi_stmt_1675: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1677_wire_constant & RPIPE_noblock_obuf_3_3_1679_wire;
      req <= phi_stmt_1675_req_0 & phi_stmt_1675_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1675",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1675_ack_0,
          idata => idata,
          odata => pkt_3_e_word_1675,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1675
    phi_stmt_1680: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1682_wire_constant & RPIPE_noblock_obuf_4_3_1684_wire;
      req <= phi_stmt_1680_req_0 & phi_stmt_1680_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1680",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1680_ack_0,
          idata => idata,
          odata => pkt_4_e_word_1680,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1680
    phi_stmt_1685: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_3_1687_wire_constant & next_active_packet_1795_1688_buffered;
      req <= phi_stmt_1685_req_0 & phi_stmt_1685_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1685",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1685_ack_0,
          idata => idata,
          odata => active_packet_1685,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1685
    phi_stmt_1689: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_8_1691_wire_constant & next_active_packet_length_1840_1692_buffered;
      req <= phi_stmt_1689_req_0 & phi_stmt_1689_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1689",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1689_ack_0,
          idata => idata,
          odata => active_packet_length_1689,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1689
    phi_stmt_1693: Block -- phi operator 
      signal idata: std_logic_vector(3 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= next_priority_index_1795_1695_buffered & R_ZERO_2_1696_wire_constant;
      req <= phi_stmt_1693_req_0 & phi_stmt_1693_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1693",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 2) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1693_ack_0,
          idata => idata,
          odata => priority_index_1693,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1693
    -- flow-through select operator MUX_1702_inst
    MUX_1702_wire <= konst_1700_wire_constant when (read_from_1_1861(0) /=  '0') else konst_1701_wire_constant;
    -- flow-through select operator MUX_1706_inst
    MUX_1706_wire <= konst_1704_wire_constant when (read_from_2_1869(0) /=  '0') else konst_1705_wire_constant;
    -- flow-through select operator MUX_1711_inst
    MUX_1711_wire <= konst_1709_wire_constant when (read_from_3_1877(0) /=  '0') else konst_1710_wire_constant;
    -- flow-through select operator MUX_1715_inst
    MUX_1715_wire <= konst_1713_wire_constant when (read_from_4_1885(0) /=  '0') else konst_1714_wire_constant;
    -- flow-through select operator MUX_1763_inst
    MUX_1763_wire <= p1_valid_1729 when (EQ_u3_u1_1760_wire(0) /=  '0') else konst_1762_wire_constant;
    -- flow-through select operator MUX_1769_inst
    MUX_1769_wire <= p2_valid_1734 when (EQ_u3_u1_1766_wire(0) /=  '0') else konst_1768_wire_constant;
    -- flow-through select operator MUX_1776_inst
    MUX_1776_wire <= p3_valid_1739 when (EQ_u3_u1_1773_wire(0) /=  '0') else konst_1775_wire_constant;
    -- flow-through select operator MUX_1782_inst
    MUX_1782_wire <= p4_valid_1744 when (EQ_u3_u1_1779_wire(0) /=  '0') else konst_1781_wire_constant;
    -- flow-through select operator MUX_1813_inst
    MUX_1813_wire <= slice_1811_wire when (EQ_u3_u1_1809_wire(0) /=  '0') else konst_1812_wire_constant;
    -- flow-through select operator MUX_1820_inst
    MUX_1820_wire <= slice_1818_wire when (EQ_u3_u1_1816_wire(0) /=  '0') else konst_1819_wire_constant;
    -- flow-through select operator MUX_1828_inst
    MUX_1828_wire <= slice_1826_wire when (EQ_u3_u1_1824_wire(0) /=  '0') else konst_1827_wire_constant;
    -- flow-through select operator MUX_1835_inst
    MUX_1835_wire <= slice_1833_wire when (EQ_u3_u1_1831_wire(0) /=  '0') else konst_1834_wire_constant;
    -- flow-through select operator MUX_1839_inst
    next_active_packet_length_1840 <= OR_u8_u8_1837_wire when (started_new_packet_1804(0) /=  '0') else active_packet_length_1689;
    -- flow-through select operator MUX_1851_inst
    MUX_1851_wire <= SUB_u8_u8_1849_wire when (valid_active_pkt_word_read_1785(0) /=  '0') else down_counter_1661;
    -- flow-through select operator MUX_1852_inst
    next_down_counter_1853 <= SUB_u8_u8_1845_wire when (started_new_packet_1804(0) /=  '0') else MUX_1851_wire;
    -- flow-through select operator MUX_1893_inst
    MUX_1893_wire <= slice_1891_wire when (EQ_u3_u1_1889_wire(0) /=  '0') else konst_1892_wire_constant;
    -- flow-through select operator MUX_1900_inst
    MUX_1900_wire <= slice_1898_wire when (EQ_u3_u1_1896_wire(0) /=  '0') else konst_1899_wire_constant;
    -- flow-through select operator MUX_1908_inst
    MUX_1908_wire <= slice_1906_wire when (EQ_u3_u1_1904_wire(0) /=  '0') else konst_1907_wire_constant;
    -- flow-through select operator MUX_1915_inst
    MUX_1915_wire <= slice_1913_wire when (EQ_u3_u1_1911_wire(0) /=  '0') else konst_1914_wire_constant;
    -- flow-through select operator MUX_1925_inst
    MUX_1925_wire <= p1_valid_1729 when (EQ_u3_u1_1922_wire(0) /=  '0') else konst_1924_wire_constant;
    -- flow-through select operator MUX_1931_inst
    MUX_1931_wire <= p2_valid_1734 when (EQ_u3_u1_1928_wire(0) /=  '0') else konst_1930_wire_constant;
    -- flow-through select operator MUX_1938_inst
    MUX_1938_wire <= p3_valid_1739 when (EQ_u3_u1_1935_wire(0) /=  '0') else konst_1937_wire_constant;
    -- flow-through select operator MUX_1944_inst
    MUX_1944_wire <= p4_valid_1744 when (EQ_u3_u1_1941_wire(0) /=  '0') else konst_1943_wire_constant;
    -- flow-through slice operator slice_1811_inst
    slice_1811_wire <= pkt_1_e_word_1665(15 downto 8);
    -- flow-through slice operator slice_1818_inst
    slice_1818_wire <= pkt_2_e_word_1670(15 downto 8);
    -- flow-through slice operator slice_1826_inst
    slice_1826_wire <= pkt_3_e_word_1675(15 downto 8);
    -- flow-through slice operator slice_1833_inst
    slice_1833_wire <= pkt_4_e_word_1680(15 downto 8);
    -- flow-through slice operator slice_1891_inst
    slice_1891_wire <= pkt_1_e_word_1665(31 downto 0);
    -- flow-through slice operator slice_1898_inst
    slice_1898_wire <= pkt_2_e_word_1670(31 downto 0);
    -- flow-through slice operator slice_1906_inst
    slice_1906_wire <= pkt_3_e_word_1675(31 downto 0);
    -- flow-through slice operator slice_1913_inst
    slice_1913_wire <= pkt_4_e_word_1680(31 downto 0);
    next_active_packet_1795_1688_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_active_packet_1795_1688_buf_req_0;
      next_active_packet_1795_1688_buf_ack_0<= wack(0);
      rreq(0) <= next_active_packet_1795_1688_buf_req_1;
      next_active_packet_1795_1688_buf_ack_1<= rack(0);
      next_active_packet_1795_1688_buf : InterlockBuffer generic map ( -- 
        name => "next_active_packet_1795_1688_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_active_packet_1795,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_active_packet_1795_1688_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_active_packet_length_1840_1692_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_active_packet_length_1840_1692_buf_req_0;
      next_active_packet_length_1840_1692_buf_ack_0<= wack(0);
      rreq(0) <= next_active_packet_length_1840_1692_buf_req_1;
      next_active_packet_length_1840_1692_buf_ack_1<= rack(0);
      next_active_packet_length_1840_1692_buf : InterlockBuffer generic map ( -- 
        name => "next_active_packet_length_1840_1692_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_active_packet_length_1840,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_active_packet_length_1840_1692_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_down_counter_1853_1664_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_down_counter_1853_1664_buf_req_0;
      next_down_counter_1853_1664_buf_ack_0<= wack(0);
      rreq(0) <= next_down_counter_1853_1664_buf_req_1;
      next_down_counter_1853_1664_buf_ack_1<= rack(0);
      next_down_counter_1853_1664_buf : InterlockBuffer generic map ( -- 
        name => "next_down_counter_1853_1664_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_down_counter_1853,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_down_counter_1853_1664_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_priority_index_1795_1695_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_priority_index_1795_1695_buf_req_0;
      next_priority_index_1795_1695_buf_ack_0<= wack(0);
      rreq(0) <= next_priority_index_1795_1695_buf_req_1;
      next_priority_index_1795_1695_buf_ack_1<= rack(0);
      next_priority_index_1795_1695_buf : InterlockBuffer generic map ( -- 
        name => "next_priority_index_1795_1695_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 2,
        out_data_width => 2,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_priority_index_1795,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_priority_index_1795_1695_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1659_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1962_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1659_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1659_branch_req_0,
          ack0 => do_while_stmt_1659_branch_ack_0,
          ack1 => do_while_stmt_1659_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- flow through binary operator AND_u1_u1_1803_inst
    started_new_packet_1804 <= (NEQ_u3_u1_1799_wire and EQ_u8_u1_1802_wire);
    -- flow through binary operator BITSEL_u33_u1_1728_inst
    process(pkt_1_e_word_1665) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_1_e_word_1665, konst_1727_wire_constant, tmp_var);
      p1_valid_1729 <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u33_u1_1733_inst
    process(pkt_2_e_word_1670) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_2_e_word_1670, konst_1732_wire_constant, tmp_var);
      p2_valid_1734 <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u33_u1_1738_inst
    process(pkt_3_e_word_1675) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_3_e_word_1675, konst_1737_wire_constant, tmp_var);
      p3_valid_1739 <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u33_u1_1743_inst
    process(pkt_4_e_word_1680) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_4_e_word_1680, konst_1742_wire_constant, tmp_var);
      p4_valid_1744 <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1760_inst
    process(active_packet_1685) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1685, konst_1759_wire_constant, tmp_var);
      EQ_u3_u1_1760_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1766_inst
    process(active_packet_1685) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1685, konst_1765_wire_constant, tmp_var);
      EQ_u3_u1_1766_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1773_inst
    process(active_packet_1685) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1685, konst_1772_wire_constant, tmp_var);
      EQ_u3_u1_1773_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1779_inst
    process(active_packet_1685) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1685, konst_1778_wire_constant, tmp_var);
      EQ_u3_u1_1779_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1809_inst
    process(next_active_packet_1795) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1795, konst_1808_wire_constant, tmp_var);
      EQ_u3_u1_1809_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1816_inst
    process(next_active_packet_1795) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1795, konst_1815_wire_constant, tmp_var);
      EQ_u3_u1_1816_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1824_inst
    process(next_active_packet_1795) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1795, konst_1823_wire_constant, tmp_var);
      EQ_u3_u1_1824_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1831_inst
    process(next_active_packet_1795) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1795, konst_1830_wire_constant, tmp_var);
      EQ_u3_u1_1831_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1859_inst
    process(next_active_packet_1795) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1795, konst_1858_wire_constant, tmp_var);
      EQ_u3_u1_1859_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1867_inst
    process(next_active_packet_1795) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1795, konst_1866_wire_constant, tmp_var);
      EQ_u3_u1_1867_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1875_inst
    process(next_active_packet_1795) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1795, konst_1874_wire_constant, tmp_var);
      EQ_u3_u1_1875_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1883_inst
    process(next_active_packet_1795) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1795, konst_1882_wire_constant, tmp_var);
      EQ_u3_u1_1883_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1889_inst
    process(next_active_packet_1795) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1795, konst_1888_wire_constant, tmp_var);
      EQ_u3_u1_1889_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1896_inst
    process(next_active_packet_1795) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1795, konst_1895_wire_constant, tmp_var);
      EQ_u3_u1_1896_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1904_inst
    process(next_active_packet_1795) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1795, konst_1903_wire_constant, tmp_var);
      EQ_u3_u1_1904_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1911_inst
    process(next_active_packet_1795) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1795, konst_1910_wire_constant, tmp_var);
      EQ_u3_u1_1911_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1922_inst
    process(next_active_packet_1795) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1795, konst_1921_wire_constant, tmp_var);
      EQ_u3_u1_1922_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1928_inst
    process(next_active_packet_1795) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1795, konst_1927_wire_constant, tmp_var);
      EQ_u3_u1_1928_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1935_inst
    process(next_active_packet_1795) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1795, konst_1934_wire_constant, tmp_var);
      EQ_u3_u1_1935_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_1941_inst
    process(next_active_packet_1795) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1795, konst_1940_wire_constant, tmp_var);
      EQ_u3_u1_1941_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u8_u1_1802_inst
    process(down_counter_1661) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(down_counter_1661, konst_1801_wire_constant, tmp_var);
      EQ_u8_u1_1802_wire <= tmp_var; --
    end process;
    -- flow through binary operator NEQ_u3_u1_1799_inst
    process(next_active_packet_1795) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(next_active_packet_1795, konst_1798_wire_constant, tmp_var);
      NEQ_u3_u1_1799_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1856_inst
    process(p1_valid_1729) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p1_valid_1729, tmp_var);
      NOT_u1_u1_1856_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1864_inst
    process(p2_valid_1734) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p2_valid_1734, tmp_var);
      NOT_u1_u1_1864_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1872_inst
    process(p3_valid_1739) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p3_valid_1739, tmp_var);
      NOT_u1_u1_1872_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1880_inst
    process(p4_valid_1744) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p4_valid_1744, tmp_var);
      NOT_u1_u1_1880_wire <= tmp_var; -- 
    end process;
    -- flow through binary operator OR_u1_u1_1770_inst
    OR_u1_u1_1770_wire <= (MUX_1763_wire or MUX_1769_wire);
    -- flow through binary operator OR_u1_u1_1783_inst
    OR_u1_u1_1783_wire <= (MUX_1776_wire or MUX_1782_wire);
    -- flow through binary operator OR_u1_u1_1784_inst
    valid_active_pkt_word_read_1785 <= (OR_u1_u1_1770_wire or OR_u1_u1_1783_wire);
    -- flow through binary operator OR_u1_u1_1860_inst
    read_from_1_1861 <= (NOT_u1_u1_1856_wire or EQ_u3_u1_1859_wire);
    -- flow through binary operator OR_u1_u1_1868_inst
    read_from_2_1869 <= (NOT_u1_u1_1864_wire or EQ_u3_u1_1867_wire);
    -- flow through binary operator OR_u1_u1_1876_inst
    read_from_3_1877 <= (NOT_u1_u1_1872_wire or EQ_u3_u1_1875_wire);
    -- flow through binary operator OR_u1_u1_1884_inst
    read_from_4_1885 <= (NOT_u1_u1_1880_wire or EQ_u3_u1_1883_wire);
    -- flow through binary operator OR_u1_u1_1932_inst
    OR_u1_u1_1932_wire <= (MUX_1925_wire or MUX_1931_wire);
    -- flow through binary operator OR_u1_u1_1945_inst
    OR_u1_u1_1945_wire <= (MUX_1938_wire or MUX_1944_wire);
    -- flow through binary operator OR_u1_u1_1946_inst
    send_flag_1947 <= (OR_u1_u1_1932_wire or OR_u1_u1_1945_wire);
    -- flow through binary operator OR_u32_u32_1901_inst
    OR_u32_u32_1901_wire <= (MUX_1893_wire or MUX_1900_wire);
    -- flow through binary operator OR_u32_u32_1916_inst
    OR_u32_u32_1916_wire <= (MUX_1908_wire or MUX_1915_wire);
    -- flow through binary operator OR_u32_u32_1917_inst
    data_to_out_1918 <= (OR_u32_u32_1901_wire or OR_u32_u32_1916_wire);
    -- flow through binary operator OR_u8_u8_1707_inst
    OR_u8_u8_1707_wire <= (MUX_1702_wire or MUX_1706_wire);
    -- flow through binary operator OR_u8_u8_1716_inst
    OR_u8_u8_1716_wire <= (MUX_1711_wire or MUX_1715_wire);
    -- flow through binary operator OR_u8_u8_1717_inst
    senderPort_1718 <= (OR_u8_u8_1707_wire or OR_u8_u8_1716_wire);
    -- flow through binary operator OR_u8_u8_1821_inst
    OR_u8_u8_1821_wire <= (MUX_1813_wire or MUX_1820_wire);
    -- flow through binary operator OR_u8_u8_1836_inst
    OR_u8_u8_1836_wire <= (MUX_1828_wire or MUX_1835_wire);
    -- flow through binary operator OR_u8_u8_1837_inst
    OR_u8_u8_1837_wire <= (OR_u8_u8_1821_wire or OR_u8_u8_1836_wire);
    -- flow through binary operator SUB_u8_u8_1845_inst
    SUB_u8_u8_1845_wire <= std_logic_vector(unsigned(next_active_packet_length_1840) - unsigned(konst_1844_wire_constant));
    -- flow through binary operator SUB_u8_u8_1849_inst
    SUB_u8_u8_1849_wire <= std_logic_vector(unsigned(down_counter_1661) - unsigned(konst_1848_wire_constant));
    -- shared inport operator group (0) : RPIPE_noblock_obuf_1_3_1669_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_1_3_1669_inst_req_0;
      RPIPE_noblock_obuf_1_3_1669_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_1_3_1669_inst_req_1;
      RPIPE_noblock_obuf_1_3_1669_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_1_1861(0);
      RPIPE_noblock_obuf_1_3_1669_wire <= data_out(32 downto 0);
      noblock_obuf_1_3_read_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_3_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_3_read_0: InputPortRevised -- 
        generic map ( name => "noblock_obuf_1_3_read_0", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_1_3_pipe_read_req(0),
          oack => noblock_obuf_1_3_pipe_read_ack(0),
          odata => noblock_obuf_1_3_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_noblock_obuf_2_3_1674_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_2_3_1674_inst_req_0;
      RPIPE_noblock_obuf_2_3_1674_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_2_3_1674_inst_req_1;
      RPIPE_noblock_obuf_2_3_1674_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_2_1869(0);
      RPIPE_noblock_obuf_2_3_1674_wire <= data_out(32 downto 0);
      noblock_obuf_2_3_read_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_3_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_3_read_1: InputPortRevised -- 
        generic map ( name => "noblock_obuf_2_3_read_1", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_2_3_pipe_read_req(0),
          oack => noblock_obuf_2_3_pipe_read_ack(0),
          odata => noblock_obuf_2_3_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_noblock_obuf_3_3_1679_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_3_3_1679_inst_req_0;
      RPIPE_noblock_obuf_3_3_1679_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_3_3_1679_inst_req_1;
      RPIPE_noblock_obuf_3_3_1679_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_3_1877(0);
      RPIPE_noblock_obuf_3_3_1679_wire <= data_out(32 downto 0);
      noblock_obuf_3_3_read_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_3_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_3_read_2: InputPortRevised -- 
        generic map ( name => "noblock_obuf_3_3_read_2", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_3_3_pipe_read_req(0),
          oack => noblock_obuf_3_3_pipe_read_ack(0),
          odata => noblock_obuf_3_3_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_noblock_obuf_4_3_1684_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_4_3_1684_inst_req_0;
      RPIPE_noblock_obuf_4_3_1684_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_4_3_1684_inst_req_1;
      RPIPE_noblock_obuf_4_3_1684_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_4_1885(0);
      RPIPE_noblock_obuf_4_3_1684_wire <= data_out(32 downto 0);
      noblock_obuf_4_3_read_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_3_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_3_read_3: InputPortRevised -- 
        generic map ( name => "noblock_obuf_4_3_read_3", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_4_3_pipe_read_req(0),
          oack => noblock_obuf_4_3_pipe_read_ack(0),
          odata => noblock_obuf_4_3_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_out_data_3_1949_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_out_data_3_1949_inst_req_0;
      WPIPE_out_data_3_1949_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_out_data_3_1949_inst_req_1;
      WPIPE_out_data_3_1949_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_flag_1947(0);
      data_in <= data_to_out_1918;
      out_data_3_write_0_gI: SplitGuardInterface generic map(name => "out_data_3_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      out_data_3_write_0: OutputPortRevised -- 
        generic map ( name => "out_data_3", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => out_data_3_pipe_write_req(0),
          oack => out_data_3_pipe_write_ack(0),
          odata => out_data_3_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_1724_call 
    updateCounter_call_group_0: Block -- 
      signal data_in: std_logic_vector(16 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1724_call_req_0;
      call_stmt_1724_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1724_call_req_1;
      call_stmt_1724_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      updateCounter_call_group_0_gI: SplitGuardInterface generic map(name => "updateCounter_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= senderPort_1718 & konst_1720_wire_constant & type_cast_1722_wire_constant;
      continue_1724 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 17,
        owidth => 17,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => updateCounter_call_reqs(0),
          ackR => updateCounter_call_acks(0),
          dataR => updateCounter_call_data(16 downto 0),
          tagR => updateCounter_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => updateCounter_return_acks(0), -- cross-over
          ackL => updateCounter_return_reqs(0), -- cross-over
          dataL => updateCounter_return_data(0 downto 0),
          tagL => updateCounter_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    volatile_operator_prioritySelect_5714: prioritySelect_Volatile port map(down_counter => down_counter_1661, active_packet => active_packet_1685, priority_index => priority_index_1693, p1_valid => p1_valid_1729, p2_valid => p2_valid_1734, p3_valid => p3_valid_1739, p4_valid => p4_valid_1744, next_active_packet => next_active_packet_1795, next_priority_index => next_priority_index_1795); 
    -- 
  end Block; -- data_path
  -- 
end outputPort_3_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity outputPort_4_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    noblock_obuf_1_4_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_4_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_3_4_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_4_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_2_4_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_4_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_4_4_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_4_pipe_read_data : in   std_logic_vector(32 downto 0);
    out_data_4_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_data_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_data_4_pipe_write_data : out  std_logic_vector(31 downto 0);
    updateCounter_call_reqs : out  std_logic_vector(0 downto 0);
    updateCounter_call_acks : in   std_logic_vector(0 downto 0);
    updateCounter_call_data : out  std_logic_vector(16 downto 0);
    updateCounter_call_tag  :  out  std_logic_vector(0 downto 0);
    updateCounter_return_reqs : out  std_logic_vector(0 downto 0);
    updateCounter_return_acks : in   std_logic_vector(0 downto 0);
    updateCounter_return_data : in   std_logic_vector(0 downto 0);
    updateCounter_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity outputPort_4_Daemon;
architecture outputPort_4_Daemon_arch of outputPort_4_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal outputPort_4_Daemon_CP_3687_start: Boolean;
  signal outputPort_4_Daemon_CP_3687_symbol: Boolean;
  -- volatile/operator module components. 
  component updateCounter is -- 
    generic (tag_length : integer); 
    port ( -- 
      input_port : in  std_logic_vector(7 downto 0);
      output_port : in  std_logic_vector(7 downto 0);
      up : in  std_logic_vector(0 downto 0);
      continue : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(3 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(1 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(1 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component prioritySelect_Volatile is -- 
    port ( -- 
      down_counter : in  std_logic_vector(7 downto 0);
      active_packet : in  std_logic_vector(2 downto 0);
      priority_index : in  std_logic_vector(1 downto 0);
      p1_valid : in  std_logic_vector(0 downto 0);
      p2_valid : in  std_logic_vector(0 downto 0);
      p3_valid : in  std_logic_vector(0 downto 0);
      p4_valid : in  std_logic_vector(0 downto 0);
      next_active_packet : out  std_logic_vector(2 downto 0);
      next_priority_index : out  std_logic_vector(1 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal next_priority_index_2103_2004_buf_ack_0 : boolean;
  signal do_while_stmt_1967_branch_req_0 : boolean;
  signal next_priority_index_2103_2004_buf_ack_1 : boolean;
  signal next_priority_index_2103_2004_buf_req_1 : boolean;
  signal call_stmt_2032_call_req_0 : boolean;
  signal phi_stmt_2001_req_0 : boolean;
  signal call_stmt_2032_call_req_1 : boolean;
  signal call_stmt_2032_call_ack_0 : boolean;
  signal phi_stmt_2001_ack_0 : boolean;
  signal next_priority_index_2103_2004_buf_req_0 : boolean;
  signal phi_stmt_2001_req_1 : boolean;
  signal phi_stmt_1969_req_1 : boolean;
  signal phi_stmt_1969_ack_0 : boolean;
  signal next_down_counter_2161_1972_buf_req_1 : boolean;
  signal next_down_counter_2161_1972_buf_ack_1 : boolean;
  signal phi_stmt_1969_req_0 : boolean;
  signal next_down_counter_2161_1972_buf_req_0 : boolean;
  signal next_down_counter_2161_1972_buf_ack_0 : boolean;
  signal phi_stmt_1973_req_1 : boolean;
  signal phi_stmt_1973_req_0 : boolean;
  signal phi_stmt_1973_ack_0 : boolean;
  signal phi_stmt_1983_ack_0 : boolean;
  signal RPIPE_noblock_obuf_1_4_1977_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_1_4_1977_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_1_4_1977_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_1_4_1977_inst_ack_1 : boolean;
  signal phi_stmt_1978_req_1 : boolean;
  signal phi_stmt_1978_req_0 : boolean;
  signal phi_stmt_1978_ack_0 : boolean;
  signal do_while_stmt_1967_branch_ack_1 : boolean;
  signal do_while_stmt_1967_branch_ack_0 : boolean;
  signal WPIPE_out_data_4_2257_inst_ack_1 : boolean;
  signal WPIPE_out_data_4_2257_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_2_4_1982_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_2_4_1982_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_2_4_1982_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_2_4_1982_inst_ack_1 : boolean;
  signal WPIPE_out_data_4_2257_inst_ack_0 : boolean;
  signal WPIPE_out_data_4_2257_inst_req_0 : boolean;
  signal phi_stmt_1983_req_1 : boolean;
  signal phi_stmt_1983_req_0 : boolean;
  signal call_stmt_2032_call_ack_1 : boolean;
  signal RPIPE_noblock_obuf_3_4_1987_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_3_4_1987_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_3_4_1987_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_3_4_1987_inst_ack_1 : boolean;
  signal phi_stmt_1988_req_1 : boolean;
  signal phi_stmt_1988_req_0 : boolean;
  signal phi_stmt_1988_ack_0 : boolean;
  signal RPIPE_noblock_obuf_4_4_1992_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_4_4_1992_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_4_4_1992_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_4_4_1992_inst_ack_1 : boolean;
  signal phi_stmt_1993_req_1 : boolean;
  signal phi_stmt_1993_req_0 : boolean;
  signal phi_stmt_1993_ack_0 : boolean;
  signal next_active_packet_2103_1996_buf_req_0 : boolean;
  signal next_active_packet_2103_1996_buf_ack_0 : boolean;
  signal next_active_packet_2103_1996_buf_req_1 : boolean;
  signal next_active_packet_2103_1996_buf_ack_1 : boolean;
  signal phi_stmt_1997_req_1 : boolean;
  signal phi_stmt_1997_req_0 : boolean;
  signal phi_stmt_1997_ack_0 : boolean;
  signal next_active_packet_length_2148_2000_buf_req_0 : boolean;
  signal next_active_packet_length_2148_2000_buf_ack_0 : boolean;
  signal next_active_packet_length_2148_2000_buf_req_1 : boolean;
  signal next_active_packet_length_2148_2000_buf_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "outputPort_4_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  outputPort_4_Daemon_CP_3687_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "outputPort_4_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_4_Daemon_CP_3687_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= outputPort_4_Daemon_CP_3687_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_4_Daemon_CP_3687_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  outputPort_4_Daemon_CP_3687: Block -- control-path 
    signal outputPort_4_Daemon_CP_3687_elements: BooleanArray(185 downto 0);
    -- 
  begin -- 
    outputPort_4_Daemon_CP_3687_elements(0) <= outputPort_4_Daemon_CP_3687_start;
    outputPort_4_Daemon_CP_3687_symbol <= outputPort_4_Daemon_CP_3687_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1966/branch_block_stmt_1966__entry__
      -- CP-element group 0: 	 branch_block_stmt_1966/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1966/do_while_stmt_1967__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	185 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_1966/$exit
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1966/do_while_stmt_1967__exit__
      -- CP-element group 1: 	 branch_block_stmt_1966/branch_block_stmt_1966__exit__
      -- 
    outputPort_4_Daemon_CP_3687_elements(1) <= outputPort_4_Daemon_CP_3687_elements(185);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967__entry__
      -- CP-element group 2: 	 branch_block_stmt_1966/do_while_stmt_1967/$entry
      -- 
    outputPort_4_Daemon_CP_3687_elements(2) <= outputPort_4_Daemon_CP_3687_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	185 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967__exit__
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1966/do_while_stmt_1967/loop_back
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	183 
    -- CP-element group 5: 	184 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1966/do_while_stmt_1967/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1966/do_while_stmt_1967/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_1966/do_while_stmt_1967/loop_exit/$entry
      -- 
    outputPort_4_Daemon_CP_3687_elements(5) <= outputPort_4_Daemon_CP_3687_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	182 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1966/do_while_stmt_1967/loop_body_done
      -- 
    outputPort_4_Daemon_CP_3687_elements(6) <= outputPort_4_Daemon_CP_3687_elements(182);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	143 
    -- CP-element group 7: 	161 
    -- CP-element group 7: 	125 
    -- CP-element group 7: 	22 
    -- CP-element group 7: 	41 
    -- CP-element group 7: 	62 
    -- CP-element group 7: 	83 
    -- CP-element group 7: 	104 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/back_edge_to_loop_body
      -- 
    outputPort_4_Daemon_CP_3687_elements(7) <= outputPort_4_Daemon_CP_3687_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	127 
    -- CP-element group 8: 	163 
    -- CP-element group 8: 	145 
    -- CP-element group 8: 	24 
    -- CP-element group 8: 	43 
    -- CP-element group 8: 	64 
    -- CP-element group 8: 	85 
    -- CP-element group 8: 	106 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/first_time_through_loop_body
      -- 
    outputPort_4_Daemon_CP_3687_elements(8) <= outputPort_4_Daemon_CP_3687_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	119 
    -- CP-element group 9: 	156 
    -- CP-element group 9: 	157 
    -- CP-element group 9: 	139 
    -- CP-element group 9: 	120 
    -- CP-element group 9: 	181 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	17 
    -- CP-element group 9: 	35 
    -- CP-element group 9: 	36 
    -- CP-element group 9: 	138 
    -- CP-element group 9: 	56 
    -- CP-element group 9: 	57 
    -- CP-element group 9: 	77 
    -- CP-element group 9: 	78 
    -- CP-element group 9: 	98 
    -- CP-element group 9: 	99 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/$entry
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	181 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/condition_evaluated
      -- 
    condition_evaluated_3711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(10), ack => do_while_stmt_1967_branch_req_0); -- 
    outputPort_4_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(181) & outputPort_4_Daemon_CP_3687_elements(15);
      gj_outputPort_4_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	119 
    -- CP-element group 11: 	156 
    -- CP-element group 11: 	16 
    -- CP-element group 11: 	35 
    -- CP-element group 11: 	138 
    -- CP-element group 11: 	56 
    -- CP-element group 11: 	77 
    -- CP-element group 11: 	98 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	121 
    -- CP-element group 11: 	140 
    -- CP-element group 11: 	18 
    -- CP-element group 11: 	37 
    -- CP-element group 11: 	58 
    -- CP-element group 11: 	79 
    -- CP-element group 11: 	100 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_2001_sample_start__ps
      -- CP-element group 11: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/aggregated_phi_sample_req
      -- 
    outputPort_4_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 1);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(119) & outputPort_4_Daemon_CP_3687_elements(156) & outputPort_4_Daemon_CP_3687_elements(16) & outputPort_4_Daemon_CP_3687_elements(35) & outputPort_4_Daemon_CP_3687_elements(138) & outputPort_4_Daemon_CP_3687_elements(56) & outputPort_4_Daemon_CP_3687_elements(77) & outputPort_4_Daemon_CP_3687_elements(98) & outputPort_4_Daemon_CP_3687_elements(15);
      gj_outputPort_4_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	141 
    -- CP-element group 12: 	158 
    -- CP-element group 12: 	122 
    -- CP-element group 12: 	19 
    -- CP-element group 12: 	38 
    -- CP-element group 12: 	59 
    -- CP-element group 12: 	80 
    -- CP-element group 12: 	101 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	182 
    -- CP-element group 12: 	13 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	119 
    -- CP-element group 12: 	156 
    -- CP-element group 12: 	16 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	138 
    -- CP-element group 12: 	56 
    -- CP-element group 12: 	77 
    -- CP-element group 12: 	98 
    -- CP-element group 12:  members (9) 
      -- CP-element group 12: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1973_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1969_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1978_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1983_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1988_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1993_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1997_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_2001_sample_completed_
      -- 
    outputPort_4_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(141) & outputPort_4_Daemon_CP_3687_elements(158) & outputPort_4_Daemon_CP_3687_elements(122) & outputPort_4_Daemon_CP_3687_elements(19) & outputPort_4_Daemon_CP_3687_elements(38) & outputPort_4_Daemon_CP_3687_elements(59) & outputPort_4_Daemon_CP_3687_elements(80) & outputPort_4_Daemon_CP_3687_elements(101);
      gj_outputPort_4_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	182 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/aggregated_phi_sample_ack_d
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(13) is a control-delay.
    cp_element_13_delay: control_delay_element  generic map(name => " 13_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_3687_elements(12), ack => outputPort_4_Daemon_CP_3687_elements(13), clk => clk, reset =>reset);
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	157 
    -- CP-element group 14: 	139 
    -- CP-element group 14: 	120 
    -- CP-element group 14: 	17 
    -- CP-element group 14: 	36 
    -- CP-element group 14: 	57 
    -- CP-element group 14: 	78 
    -- CP-element group 14: 	99 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	123 
    -- CP-element group 14: 	159 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	39 
    -- CP-element group 14: 	60 
    -- CP-element group 14: 	81 
    -- CP-element group 14: 	102 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/aggregated_phi_update_req
      -- CP-element group 14: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1997_update_start__ps
      -- 
    outputPort_4_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(157) & outputPort_4_Daemon_CP_3687_elements(139) & outputPort_4_Daemon_CP_3687_elements(120) & outputPort_4_Daemon_CP_3687_elements(17) & outputPort_4_Daemon_CP_3687_elements(36) & outputPort_4_Daemon_CP_3687_elements(57) & outputPort_4_Daemon_CP_3687_elements(78) & outputPort_4_Daemon_CP_3687_elements(99);
      gj_outputPort_4_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	124 
    -- CP-element group 15: 	142 
    -- CP-element group 15: 	160 
    -- CP-element group 15: 	21 
    -- CP-element group 15: 	40 
    -- CP-element group 15: 	61 
    -- CP-element group 15: 	82 
    -- CP-element group 15: 	103 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/aggregated_phi_update_ack
      -- 
    outputPort_4_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 7);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(124) & outputPort_4_Daemon_CP_3687_elements(142) & outputPort_4_Daemon_CP_3687_elements(160) & outputPort_4_Daemon_CP_3687_elements(21) & outputPort_4_Daemon_CP_3687_elements(40) & outputPort_4_Daemon_CP_3687_elements(61) & outputPort_4_Daemon_CP_3687_elements(82) & outputPort_4_Daemon_CP_3687_elements(103);
      gj_outputPort_4_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	11 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1969_sample_start_
      -- 
    outputPort_4_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(9) & outputPort_4_Daemon_CP_3687_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	9 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	176 
    -- CP-element group 17: 	179 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	14 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1969_update_start_
      -- 
    outputPort_4_Daemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(9) & outputPort_4_Daemon_CP_3687_elements(176) & outputPort_4_Daemon_CP_3687_elements(179);
      gj_outputPort_4_Daemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	11 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1969_sample_start__ps
      -- 
    outputPort_4_Daemon_CP_3687_elements(18) <= outputPort_4_Daemon_CP_3687_elements(11);
    -- CP-element group 19:  join  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	12 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1969_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(19) is bound as output of CP function.
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	14 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1969_update_start__ps
      -- 
    outputPort_4_Daemon_CP_3687_elements(20) <= outputPort_4_Daemon_CP_3687_elements(14);
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	174 
    -- CP-element group 21: 	178 
    -- CP-element group 21: 	15 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1969_update_completed__ps
      -- CP-element group 21: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1969_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(21) is bound as output of CP function.
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	7 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1969_loopback_trigger
      -- 
    outputPort_4_Daemon_CP_3687_elements(22) <= outputPort_4_Daemon_CP_3687_elements(7);
    -- CP-element group 23:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1969_loopback_sample_req_ps
      -- CP-element group 23: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1969_loopback_sample_req
      -- 
    phi_stmt_1969_loopback_sample_req_3727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1969_loopback_sample_req_3727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(23), ack => phi_stmt_1969_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(23) is bound as output of CP function.
    -- CP-element group 24:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	8 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1969_entry_trigger
      -- 
    outputPort_4_Daemon_CP_3687_elements(24) <= outputPort_4_Daemon_CP_3687_elements(8);
    -- CP-element group 25:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1969_entry_sample_req_ps
      -- CP-element group 25: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1969_entry_sample_req
      -- 
    phi_stmt_1969_entry_sample_req_3730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1969_entry_sample_req_3730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(25), ack => phi_stmt_1969_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1969_phi_mux_ack_ps
      -- CP-element group 26: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1969_phi_mux_ack
      -- 
    phi_stmt_1969_phi_mux_ack_3733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1969_ack_0, ack => outputPort_4_Daemon_CP_3687_elements(26)); -- 
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_8_1971_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_8_1971_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_8_1971_sample_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_8_1971_sample_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_8_1971_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_8_1971_update_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	30 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_8_1971_update_completed__ps
      -- 
    outputPort_4_Daemon_CP_3687_elements(29) <= outputPort_4_Daemon_CP_3687_elements(30);
    -- CP-element group 30:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	29 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_8_1971_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(30) is a control-delay.
    cp_element_30_delay: control_delay_element  generic map(name => " 30_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_3687_elements(28), ack => outputPort_4_Daemon_CP_3687_elements(30), clk => clk, reset =>reset);
    -- CP-element group 31:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_down_counter_1972_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_down_counter_1972_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_down_counter_1972_sample_start__ps
      -- CP-element group 31: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_down_counter_1972_Sample/req
      -- 
    req_3754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(31), ack => next_down_counter_2161_1972_buf_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_down_counter_1972_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_down_counter_1972_update_start__ps
      -- CP-element group 32: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_down_counter_1972_Update/req
      -- CP-element group 32: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_down_counter_1972_Update/$entry
      -- 
    req_3759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(32), ack => next_down_counter_2161_1972_buf_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_down_counter_1972_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_down_counter_1972_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_down_counter_1972_sample_completed__ps
      -- CP-element group 33: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_down_counter_1972_Sample/ack
      -- 
    ack_3755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_2161_1972_buf_ack_0, ack => outputPort_4_Daemon_CP_3687_elements(33)); -- 
    -- CP-element group 34:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_down_counter_1972_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_down_counter_1972_update_completed__ps
      -- CP-element group 34: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_down_counter_1972_Update/ack
      -- CP-element group 34: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_down_counter_1972_Update/$exit
      -- 
    ack_3760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_2161_1972_buf_ack_1, ack => outputPort_4_Daemon_CP_3687_elements(34)); -- 
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	12 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	11 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1973_sample_start_
      -- 
    outputPort_4_Daemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(9) & outputPort_4_Daemon_CP_3687_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	9 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	176 
    -- CP-element group 36: 	179 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	14 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1973_update_start_
      -- 
    outputPort_4_Daemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(9) & outputPort_4_Daemon_CP_3687_elements(176) & outputPort_4_Daemon_CP_3687_elements(179);
      gj_outputPort_4_Daemon_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	11 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1973_sample_start__ps
      -- 
    outputPort_4_Daemon_CP_3687_elements(37) <= outputPort_4_Daemon_CP_3687_elements(11);
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	12 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1973_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(38) is bound as output of CP function.
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	14 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1973_update_start__ps
      -- 
    outputPort_4_Daemon_CP_3687_elements(39) <= outputPort_4_Daemon_CP_3687_elements(14);
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	174 
    -- CP-element group 40: 	178 
    -- CP-element group 40: 	15 
    -- CP-element group 40:  members (2) 
      -- CP-element group 40: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1973_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1973_update_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(40) is bound as output of CP function.
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	7 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1973_loopback_trigger
      -- 
    outputPort_4_Daemon_CP_3687_elements(41) <= outputPort_4_Daemon_CP_3687_elements(7);
    -- CP-element group 42:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1973_loopback_sample_req
      -- CP-element group 42: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1973_loopback_sample_req_ps
      -- 
    phi_stmt_1973_loopback_sample_req_3771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1973_loopback_sample_req_3771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(42), ack => phi_stmt_1973_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(42) is bound as output of CP function.
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	8 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1973_entry_trigger
      -- 
    outputPort_4_Daemon_CP_3687_elements(43) <= outputPort_4_Daemon_CP_3687_elements(8);
    -- CP-element group 44:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1973_entry_sample_req
      -- CP-element group 44: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1973_entry_sample_req_ps
      -- 
    phi_stmt_1973_entry_sample_req_3774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1973_entry_sample_req_3774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(44), ack => phi_stmt_1973_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(44) is bound as output of CP function.
    -- CP-element group 45:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1973_phi_mux_ack
      -- CP-element group 45: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1973_phi_mux_ack_ps
      -- 
    phi_stmt_1973_phi_mux_ack_3777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1973_ack_0, ack => outputPort_4_Daemon_CP_3687_elements(45)); -- 
    -- CP-element group 46:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (4) 
      -- CP-element group 46: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1975_sample_start__ps
      -- CP-element group 46: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1975_sample_completed__ps
      -- CP-element group 46: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1975_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1975_sample_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1975_update_start__ps
      -- CP-element group 47: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1975_update_start_
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	49 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1975_update_completed__ps
      -- 
    outputPort_4_Daemon_CP_3687_elements(48) <= outputPort_4_Daemon_CP_3687_elements(49);
    -- CP-element group 49:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	48 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1975_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(49) is a control-delay.
    cp_element_49_delay: control_delay_element  generic map(name => " 49_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_3687_elements(47), ack => outputPort_4_Daemon_CP_3687_elements(49), clk => clk, reset =>reset);
    -- CP-element group 50:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_1_4_1977_sample_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_1_4_1977_update_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(51) is bound as output of CP function.
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	55 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_1_4_1977_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_1_4_1977_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_1_4_1977_Sample/rr
      -- 
    rr_3798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(52), ack => RPIPE_noblock_obuf_1_4_1977_inst_req_0); -- 
    outputPort_4_Daemon_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(50) & outputPort_4_Daemon_CP_3687_elements(55);
      gj_outputPort_4_Daemon_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: 	54 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_1_4_1977_update_start_
      -- CP-element group 53: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_1_4_1977_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_1_4_1977_Update/cr
      -- 
    cr_3803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(53), ack => RPIPE_noblock_obuf_1_4_1977_inst_req_1); -- 
    outputPort_4_Daemon_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(51) & outputPort_4_Daemon_CP_3687_elements(54);
      gj_outputPort_4_Daemon_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	53 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_1_4_1977_sample_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_1_4_1977_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_1_4_1977_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_1_4_1977_Sample/ra
      -- 
    ra_3799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_4_1977_inst_ack_0, ack => outputPort_4_Daemon_CP_3687_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: marked-successors 
    -- CP-element group 55: 	52 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_1_4_1977_update_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_1_4_1977_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_1_4_1977_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_1_4_1977_Update/ca
      -- 
    ca_3804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_4_1977_inst_ack_1, ack => outputPort_4_Daemon_CP_3687_elements(55)); -- 
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	9 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	12 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	11 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1978_sample_start_
      -- 
    outputPort_4_Daemon_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(9) & outputPort_4_Daemon_CP_3687_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  join  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	9 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	176 
    -- CP-element group 57: 	179 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	14 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1978_update_start_
      -- 
    outputPort_4_Daemon_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(9) & outputPort_4_Daemon_CP_3687_elements(176) & outputPort_4_Daemon_CP_3687_elements(179);
      gj_outputPort_4_Daemon_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	11 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1978_sample_start__ps
      -- 
    outputPort_4_Daemon_CP_3687_elements(58) <= outputPort_4_Daemon_CP_3687_elements(11);
    -- CP-element group 59:  join  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	12 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1978_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(59) is bound as output of CP function.
    -- CP-element group 60:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	14 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1978_update_start__ps
      -- 
    outputPort_4_Daemon_CP_3687_elements(60) <= outputPort_4_Daemon_CP_3687_elements(14);
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	174 
    -- CP-element group 61: 	178 
    -- CP-element group 61: 	15 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1978_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1978_update_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(61) is bound as output of CP function.
    -- CP-element group 62:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	7 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1978_loopback_trigger
      -- 
    outputPort_4_Daemon_CP_3687_elements(62) <= outputPort_4_Daemon_CP_3687_elements(7);
    -- CP-element group 63:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1978_loopback_sample_req
      -- CP-element group 63: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1978_loopback_sample_req_ps
      -- 
    phi_stmt_1978_loopback_sample_req_3815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1978_loopback_sample_req_3815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(63), ack => phi_stmt_1978_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(63) is bound as output of CP function.
    -- CP-element group 64:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	8 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1978_entry_trigger
      -- 
    outputPort_4_Daemon_CP_3687_elements(64) <= outputPort_4_Daemon_CP_3687_elements(8);
    -- CP-element group 65:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1978_entry_sample_req
      -- CP-element group 65: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1978_entry_sample_req_ps
      -- 
    phi_stmt_1978_entry_sample_req_3818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1978_entry_sample_req_3818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(65), ack => phi_stmt_1978_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(65) is bound as output of CP function.
    -- CP-element group 66:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1978_phi_mux_ack
      -- CP-element group 66: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1978_phi_mux_ack_ps
      -- 
    phi_stmt_1978_phi_mux_ack_3821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1978_ack_0, ack => outputPort_4_Daemon_CP_3687_elements(66)); -- 
    -- CP-element group 67:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1980_sample_start__ps
      -- CP-element group 67: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1980_sample_completed__ps
      -- CP-element group 67: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1980_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1980_sample_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1980_update_start__ps
      -- CP-element group 68: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1980_update_start_
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	70 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1980_update_completed__ps
      -- 
    outputPort_4_Daemon_CP_3687_elements(69) <= outputPort_4_Daemon_CP_3687_elements(70);
    -- CP-element group 70:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	69 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1980_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(70) is a control-delay.
    cp_element_70_delay: control_delay_element  generic map(name => " 70_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_3687_elements(68), ack => outputPort_4_Daemon_CP_3687_elements(70), clk => clk, reset =>reset);
    -- CP-element group 71:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_2_4_1982_sample_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(71) is bound as output of CP function.
    -- CP-element group 72:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_2_4_1982_update_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(72) is bound as output of CP function.
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: marked-predecessors 
    -- CP-element group 73: 	76 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_2_4_1982_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_2_4_1982_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_2_4_1982_Sample/rr
      -- 
    rr_3842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(73), ack => RPIPE_noblock_obuf_2_4_1982_inst_req_0); -- 
    outputPort_4_Daemon_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(71) & outputPort_4_Daemon_CP_3687_elements(76);
      gj_outputPort_4_Daemon_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: 	75 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_2_4_1982_update_start_
      -- CP-element group 74: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_2_4_1982_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_2_4_1982_Update/cr
      -- 
    cr_3847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(74), ack => RPIPE_noblock_obuf_2_4_1982_inst_req_1); -- 
    outputPort_4_Daemon_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(72) & outputPort_4_Daemon_CP_3687_elements(75);
      gj_outputPort_4_Daemon_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	74 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_2_4_1982_sample_completed__ps
      -- CP-element group 75: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_2_4_1982_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_2_4_1982_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_2_4_1982_Sample/ra
      -- 
    ra_3843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_4_1982_inst_ack_0, ack => outputPort_4_Daemon_CP_3687_elements(75)); -- 
    -- CP-element group 76:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: marked-successors 
    -- CP-element group 76: 	73 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_2_4_1982_update_completed__ps
      -- CP-element group 76: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_2_4_1982_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_2_4_1982_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_2_4_1982_Update/ca
      -- 
    ca_3848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_4_1982_inst_ack_1, ack => outputPort_4_Daemon_CP_3687_elements(76)); -- 
    -- CP-element group 77:  join  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	9 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	12 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	11 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1983_sample_start_
      -- 
    outputPort_4_Daemon_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(9) & outputPort_4_Daemon_CP_3687_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  join  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	9 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	176 
    -- CP-element group 78: 	179 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	14 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1983_update_start_
      -- 
    outputPort_4_Daemon_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(9) & outputPort_4_Daemon_CP_3687_elements(176) & outputPort_4_Daemon_CP_3687_elements(179);
      gj_outputPort_4_Daemon_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	11 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1983_sample_start__ps
      -- 
    outputPort_4_Daemon_CP_3687_elements(79) <= outputPort_4_Daemon_CP_3687_elements(11);
    -- CP-element group 80:  join  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	12 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1983_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(80) is bound as output of CP function.
    -- CP-element group 81:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	14 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1983_update_start__ps
      -- 
    outputPort_4_Daemon_CP_3687_elements(81) <= outputPort_4_Daemon_CP_3687_elements(14);
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	174 
    -- CP-element group 82: 	178 
    -- CP-element group 82: 	15 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1983_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1983_update_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(82) is bound as output of CP function.
    -- CP-element group 83:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	7 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1983_loopback_trigger
      -- 
    outputPort_4_Daemon_CP_3687_elements(83) <= outputPort_4_Daemon_CP_3687_elements(7);
    -- CP-element group 84:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1983_loopback_sample_req
      -- CP-element group 84: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1983_loopback_sample_req_ps
      -- 
    phi_stmt_1983_loopback_sample_req_3859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1983_loopback_sample_req_3859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(84), ack => phi_stmt_1983_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(84) is bound as output of CP function.
    -- CP-element group 85:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	8 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1983_entry_trigger
      -- 
    outputPort_4_Daemon_CP_3687_elements(85) <= outputPort_4_Daemon_CP_3687_elements(8);
    -- CP-element group 86:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1983_entry_sample_req
      -- CP-element group 86: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1983_entry_sample_req_ps
      -- 
    phi_stmt_1983_entry_sample_req_3862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1983_entry_sample_req_3862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(86), ack => phi_stmt_1983_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(86) is bound as output of CP function.
    -- CP-element group 87:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1983_phi_mux_ack
      -- CP-element group 87: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1983_phi_mux_ack_ps
      -- 
    phi_stmt_1983_phi_mux_ack_3865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1983_ack_0, ack => outputPort_4_Daemon_CP_3687_elements(87)); -- 
    -- CP-element group 88:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (4) 
      -- CP-element group 88: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1985_sample_start__ps
      -- CP-element group 88: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1985_sample_completed__ps
      -- CP-element group 88: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1985_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1985_sample_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1985_update_start__ps
      -- CP-element group 89: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1985_update_start_
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(89) is bound as output of CP function.
    -- CP-element group 90:  join  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	91 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1985_update_completed__ps
      -- 
    outputPort_4_Daemon_CP_3687_elements(90) <= outputPort_4_Daemon_CP_3687_elements(91);
    -- CP-element group 91:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	90 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1985_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(91) is a control-delay.
    cp_element_91_delay: control_delay_element  generic map(name => " 91_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_3687_elements(89), ack => outputPort_4_Daemon_CP_3687_elements(91), clk => clk, reset =>reset);
    -- CP-element group 92:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_3_4_1987_sample_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(92) is bound as output of CP function.
    -- CP-element group 93:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_3_4_1987_update_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(93) is bound as output of CP function.
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	97 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_3_4_1987_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_3_4_1987_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_3_4_1987_Sample/rr
      -- 
    rr_3886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(94), ack => RPIPE_noblock_obuf_3_4_1987_inst_req_0); -- 
    outputPort_4_Daemon_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(92) & outputPort_4_Daemon_CP_3687_elements(97);
      gj_outputPort_4_Daemon_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: 	96 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_3_4_1987_update_start_
      -- CP-element group 95: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_3_4_1987_Update/$entry
      -- CP-element group 95: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_3_4_1987_Update/cr
      -- 
    cr_3891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(95), ack => RPIPE_noblock_obuf_3_4_1987_inst_req_1); -- 
    outputPort_4_Daemon_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(93) & outputPort_4_Daemon_CP_3687_elements(96);
      gj_outputPort_4_Daemon_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	95 
    -- CP-element group 96:  members (4) 
      -- CP-element group 96: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_3_4_1987_sample_completed__ps
      -- CP-element group 96: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_3_4_1987_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_3_4_1987_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_3_4_1987_Sample/ra
      -- 
    ra_3887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_4_1987_inst_ack_0, ack => outputPort_4_Daemon_CP_3687_elements(96)); -- 
    -- CP-element group 97:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: marked-successors 
    -- CP-element group 97: 	94 
    -- CP-element group 97:  members (4) 
      -- CP-element group 97: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_3_4_1987_update_completed__ps
      -- CP-element group 97: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_3_4_1987_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_3_4_1987_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_3_4_1987_Update/ca
      -- 
    ca_3892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_4_1987_inst_ack_1, ack => outputPort_4_Daemon_CP_3687_elements(97)); -- 
    -- CP-element group 98:  join  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	9 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	12 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	11 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1988_sample_start_
      -- 
    outputPort_4_Daemon_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(9) & outputPort_4_Daemon_CP_3687_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  join  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	9 
    -- CP-element group 99: marked-predecessors 
    -- CP-element group 99: 	176 
    -- CP-element group 99: 	179 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	14 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1988_update_start_
      -- 
    outputPort_4_Daemon_cp_element_group_99: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_99"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(9) & outputPort_4_Daemon_CP_3687_elements(176) & outputPort_4_Daemon_CP_3687_elements(179);
      gj_outputPort_4_Daemon_cp_element_group_99 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(99), clk => clk, reset => reset); --
    end block;
    -- CP-element group 100:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	11 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1988_sample_start__ps
      -- 
    outputPort_4_Daemon_CP_3687_elements(100) <= outputPort_4_Daemon_CP_3687_elements(11);
    -- CP-element group 101:  join  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	12 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1988_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(101) is bound as output of CP function.
    -- CP-element group 102:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	14 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1988_update_start__ps
      -- 
    outputPort_4_Daemon_CP_3687_elements(102) <= outputPort_4_Daemon_CP_3687_elements(14);
    -- CP-element group 103:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	174 
    -- CP-element group 103: 	178 
    -- CP-element group 103: 	15 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1988_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1988_update_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(103) is bound as output of CP function.
    -- CP-element group 104:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	7 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1988_loopback_trigger
      -- 
    outputPort_4_Daemon_CP_3687_elements(104) <= outputPort_4_Daemon_CP_3687_elements(7);
    -- CP-element group 105:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1988_loopback_sample_req
      -- CP-element group 105: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1988_loopback_sample_req_ps
      -- 
    phi_stmt_1988_loopback_sample_req_3903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1988_loopback_sample_req_3903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(105), ack => phi_stmt_1988_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(105) is bound as output of CP function.
    -- CP-element group 106:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	8 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1988_entry_trigger
      -- 
    outputPort_4_Daemon_CP_3687_elements(106) <= outputPort_4_Daemon_CP_3687_elements(8);
    -- CP-element group 107:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1988_entry_sample_req
      -- CP-element group 107: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1988_entry_sample_req_ps
      -- 
    phi_stmt_1988_entry_sample_req_3906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1988_entry_sample_req_3906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(107), ack => phi_stmt_1988_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(107) is bound as output of CP function.
    -- CP-element group 108:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1988_phi_mux_ack
      -- CP-element group 108: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1988_phi_mux_ack_ps
      -- 
    phi_stmt_1988_phi_mux_ack_3909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1988_ack_0, ack => outputPort_4_Daemon_CP_3687_elements(108)); -- 
    -- CP-element group 109:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (4) 
      -- CP-element group 109: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1990_sample_start__ps
      -- CP-element group 109: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1990_sample_completed__ps
      -- CP-element group 109: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1990_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1990_sample_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(109) is bound as output of CP function.
    -- CP-element group 110:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1990_update_start__ps
      -- CP-element group 110: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1990_update_start_
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(110) is bound as output of CP function.
    -- CP-element group 111:  join  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1990_update_completed__ps
      -- 
    outputPort_4_Daemon_CP_3687_elements(111) <= outputPort_4_Daemon_CP_3687_elements(112);
    -- CP-element group 112:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	111 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_33_1990_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(112) is a control-delay.
    cp_element_112_delay: control_delay_element  generic map(name => " 112_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_3687_elements(110), ack => outputPort_4_Daemon_CP_3687_elements(112), clk => clk, reset =>reset);
    -- CP-element group 113:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_4_4_1992_sample_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(113) is bound as output of CP function.
    -- CP-element group 114:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_4_4_1992_update_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(114) is bound as output of CP function.
    -- CP-element group 115:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: marked-predecessors 
    -- CP-element group 115: 	118 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_4_4_1992_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_4_4_1992_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_4_4_1992_Sample/rr
      -- 
    rr_3930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(115), ack => RPIPE_noblock_obuf_4_4_1992_inst_req_0); -- 
    outputPort_4_Daemon_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(113) & outputPort_4_Daemon_CP_3687_elements(118);
      gj_outputPort_4_Daemon_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	117 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_4_4_1992_update_start_
      -- CP-element group 116: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_4_4_1992_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_4_4_1992_Update/cr
      -- 
    cr_3935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(116), ack => RPIPE_noblock_obuf_4_4_1992_inst_req_1); -- 
    outputPort_4_Daemon_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(117) & outputPort_4_Daemon_CP_3687_elements(114);
      gj_outputPort_4_Daemon_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	116 
    -- CP-element group 117:  members (4) 
      -- CP-element group 117: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_4_4_1992_sample_completed__ps
      -- CP-element group 117: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_4_4_1992_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_4_4_1992_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_4_4_1992_Sample/ra
      -- 
    ra_3931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_4_1992_inst_ack_0, ack => outputPort_4_Daemon_CP_3687_elements(117)); -- 
    -- CP-element group 118:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: marked-successors 
    -- CP-element group 118: 	115 
    -- CP-element group 118:  members (4) 
      -- CP-element group 118: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_4_4_1992_update_completed__ps
      -- CP-element group 118: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_4_4_1992_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_4_4_1992_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/RPIPE_noblock_obuf_4_4_1992_Update/ca
      -- 
    ca_3936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_4_1992_inst_ack_1, ack => outputPort_4_Daemon_CP_3687_elements(118)); -- 
    -- CP-element group 119:  join  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	9 
    -- CP-element group 119: marked-predecessors 
    -- CP-element group 119: 	12 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	11 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1993_sample_start_
      -- 
    outputPort_4_Daemon_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(9) & outputPort_4_Daemon_CP_3687_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  join  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	9 
    -- CP-element group 120: marked-predecessors 
    -- CP-element group 120: 	176 
    -- CP-element group 120: 	179 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	14 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1993_update_start_
      -- 
    outputPort_4_Daemon_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(9) & outputPort_4_Daemon_CP_3687_elements(176) & outputPort_4_Daemon_CP_3687_elements(179);
      gj_outputPort_4_Daemon_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	11 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1993_sample_start__ps
      -- 
    outputPort_4_Daemon_CP_3687_elements(121) <= outputPort_4_Daemon_CP_3687_elements(11);
    -- CP-element group 122:  join  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	12 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1993_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(122) is bound as output of CP function.
    -- CP-element group 123:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	14 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1993_update_start__ps
      -- 
    outputPort_4_Daemon_CP_3687_elements(123) <= outputPort_4_Daemon_CP_3687_elements(14);
    -- CP-element group 124:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	174 
    -- CP-element group 124: 	178 
    -- CP-element group 124: 	15 
    -- CP-element group 124:  members (2) 
      -- CP-element group 124: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1993_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1993_update_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(124) is bound as output of CP function.
    -- CP-element group 125:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	7 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1993_loopback_trigger
      -- 
    outputPort_4_Daemon_CP_3687_elements(125) <= outputPort_4_Daemon_CP_3687_elements(7);
    -- CP-element group 126:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1993_loopback_sample_req
      -- CP-element group 126: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1993_loopback_sample_req_ps
      -- 
    phi_stmt_1993_loopback_sample_req_3947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1993_loopback_sample_req_3947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(126), ack => phi_stmt_1993_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(126) is bound as output of CP function.
    -- CP-element group 127:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	8 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1993_entry_trigger
      -- 
    outputPort_4_Daemon_CP_3687_elements(127) <= outputPort_4_Daemon_CP_3687_elements(8);
    -- CP-element group 128:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1993_entry_sample_req
      -- CP-element group 128: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1993_entry_sample_req_ps
      -- 
    phi_stmt_1993_entry_sample_req_3950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1993_entry_sample_req_3950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(128), ack => phi_stmt_1993_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(128) is bound as output of CP function.
    -- CP-element group 129:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (2) 
      -- CP-element group 129: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1993_phi_mux_ack
      -- CP-element group 129: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1993_phi_mux_ack_ps
      -- 
    phi_stmt_1993_phi_mux_ack_3953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1993_ack_0, ack => outputPort_4_Daemon_CP_3687_elements(129)); -- 
    -- CP-element group 130:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: successors 
    -- CP-element group 130:  members (4) 
      -- CP-element group 130: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_3_1995_sample_start__ps
      -- CP-element group 130: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_3_1995_sample_completed__ps
      -- CP-element group 130: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_3_1995_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_3_1995_sample_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(130) is bound as output of CP function.
    -- CP-element group 131:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (2) 
      -- CP-element group 131: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_3_1995_update_start__ps
      -- CP-element group 131: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_3_1995_update_start_
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(131) is bound as output of CP function.
    -- CP-element group 132:  join  transition  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	133 
    -- CP-element group 132: successors 
    -- CP-element group 132:  members (1) 
      -- CP-element group 132: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_3_1995_update_completed__ps
      -- 
    outputPort_4_Daemon_CP_3687_elements(132) <= outputPort_4_Daemon_CP_3687_elements(133);
    -- CP-element group 133:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	132 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_3_1995_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(133) is a control-delay.
    cp_element_133_delay: control_delay_element  generic map(name => " 133_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_3687_elements(131), ack => outputPort_4_Daemon_CP_3687_elements(133), clk => clk, reset =>reset);
    -- CP-element group 134:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (4) 
      -- CP-element group 134: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_1996_sample_start__ps
      -- CP-element group 134: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_1996_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_1996_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_1996_Sample/req
      -- 
    req_3974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(134), ack => next_active_packet_2103_1996_buf_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(134) is bound as output of CP function.
    -- CP-element group 135:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	137 
    -- CP-element group 135:  members (4) 
      -- CP-element group 135: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_1996_update_start__ps
      -- CP-element group 135: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_1996_update_start_
      -- CP-element group 135: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_1996_Update/$entry
      -- CP-element group 135: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_1996_Update/req
      -- 
    req_3979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(135), ack => next_active_packet_2103_1996_buf_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(135) is bound as output of CP function.
    -- CP-element group 136:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (4) 
      -- CP-element group 136: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_1996_sample_completed__ps
      -- CP-element group 136: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_1996_sample_completed_
      -- CP-element group 136: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_1996_Sample/$exit
      -- CP-element group 136: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_1996_Sample/ack
      -- 
    ack_3975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_2103_1996_buf_ack_0, ack => outputPort_4_Daemon_CP_3687_elements(136)); -- 
    -- CP-element group 137:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	135 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (4) 
      -- CP-element group 137: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_1996_update_completed__ps
      -- CP-element group 137: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_1996_update_completed_
      -- CP-element group 137: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_1996_Update/$exit
      -- CP-element group 137: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_1996_Update/ack
      -- 
    ack_3980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_2103_1996_buf_ack_1, ack => outputPort_4_Daemon_CP_3687_elements(137)); -- 
    -- CP-element group 138:  join  transition  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	9 
    -- CP-element group 138: marked-predecessors 
    -- CP-element group 138: 	12 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	11 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1997_sample_start_
      -- 
    outputPort_4_Daemon_cp_element_group_138: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_138"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(9) & outputPort_4_Daemon_CP_3687_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_138 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(138), clk => clk, reset => reset); --
    end block;
    -- CP-element group 139:  join  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	9 
    -- CP-element group 139: marked-predecessors 
    -- CP-element group 139: 	142 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	14 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1997_update_start_
      -- 
    outputPort_4_Daemon_cp_element_group_139: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_139"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(9) & outputPort_4_Daemon_CP_3687_elements(142);
      gj_outputPort_4_Daemon_cp_element_group_139 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(139), clk => clk, reset => reset); --
    end block;
    -- CP-element group 140:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	11 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (1) 
      -- CP-element group 140: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1997_sample_start__ps
      -- 
    outputPort_4_Daemon_CP_3687_elements(140) <= outputPort_4_Daemon_CP_3687_elements(11);
    -- CP-element group 141:  join  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	12 
    -- CP-element group 141:  members (1) 
      -- CP-element group 141: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1997_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(141) is bound as output of CP function.
    -- CP-element group 142:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	15 
    -- CP-element group 142: marked-successors 
    -- CP-element group 142: 	139 
    -- CP-element group 142:  members (2) 
      -- CP-element group 142: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1997_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1997_update_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(142) is bound as output of CP function.
    -- CP-element group 143:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	7 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1997_loopback_trigger
      -- 
    outputPort_4_Daemon_CP_3687_elements(143) <= outputPort_4_Daemon_CP_3687_elements(7);
    -- CP-element group 144:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (2) 
      -- CP-element group 144: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1997_loopback_sample_req
      -- CP-element group 144: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1997_loopback_sample_req_ps
      -- 
    phi_stmt_1997_loopback_sample_req_3991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1997_loopback_sample_req_3991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(144), ack => phi_stmt_1997_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(144) is bound as output of CP function.
    -- CP-element group 145:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	8 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (1) 
      -- CP-element group 145: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1997_entry_trigger
      -- 
    outputPort_4_Daemon_CP_3687_elements(145) <= outputPort_4_Daemon_CP_3687_elements(8);
    -- CP-element group 146:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (2) 
      -- CP-element group 146: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1997_entry_sample_req
      -- CP-element group 146: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1997_entry_sample_req_ps
      -- 
    phi_stmt_1997_entry_sample_req_3994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1997_entry_sample_req_3994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(146), ack => phi_stmt_1997_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(146) is bound as output of CP function.
    -- CP-element group 147:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (2) 
      -- CP-element group 147: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1997_phi_mux_ack
      -- CP-element group 147: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_1997_phi_mux_ack_ps
      -- 
    phi_stmt_1997_phi_mux_ack_3997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1997_ack_0, ack => outputPort_4_Daemon_CP_3687_elements(147)); -- 
    -- CP-element group 148:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (4) 
      -- CP-element group 148: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_8_1999_sample_start__ps
      -- CP-element group 148: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_8_1999_sample_completed__ps
      -- CP-element group 148: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_8_1999_sample_start_
      -- CP-element group 148: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_8_1999_sample_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(148) is bound as output of CP function.
    -- CP-element group 149:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	151 
    -- CP-element group 149:  members (2) 
      -- CP-element group 149: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_8_1999_update_start__ps
      -- CP-element group 149: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_8_1999_update_start_
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(149) is bound as output of CP function.
    -- CP-element group 150:  join  transition  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	151 
    -- CP-element group 150: successors 
    -- CP-element group 150:  members (1) 
      -- CP-element group 150: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_8_1999_update_completed__ps
      -- 
    outputPort_4_Daemon_CP_3687_elements(150) <= outputPort_4_Daemon_CP_3687_elements(151);
    -- CP-element group 151:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	149 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	150 
    -- CP-element group 151:  members (1) 
      -- CP-element group 151: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_8_1999_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(151) is a control-delay.
    cp_element_151_delay: control_delay_element  generic map(name => " 151_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_3687_elements(149), ack => outputPort_4_Daemon_CP_3687_elements(151), clk => clk, reset =>reset);
    -- CP-element group 152:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (4) 
      -- CP-element group 152: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_length_2000_sample_start__ps
      -- CP-element group 152: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_length_2000_sample_start_
      -- CP-element group 152: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_length_2000_Sample/$entry
      -- CP-element group 152: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_length_2000_Sample/req
      -- 
    req_4018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(152), ack => next_active_packet_length_2148_2000_buf_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(152) is bound as output of CP function.
    -- CP-element group 153:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	155 
    -- CP-element group 153:  members (4) 
      -- CP-element group 153: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_length_2000_update_start__ps
      -- CP-element group 153: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_length_2000_update_start_
      -- CP-element group 153: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_length_2000_Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_length_2000_Update/req
      -- 
    req_4023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(153), ack => next_active_packet_length_2148_2000_buf_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(153) is bound as output of CP function.
    -- CP-element group 154:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	152 
    -- CP-element group 154: successors 
    -- CP-element group 154:  members (4) 
      -- CP-element group 154: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_length_2000_sample_completed__ps
      -- CP-element group 154: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_length_2000_sample_completed_
      -- CP-element group 154: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_length_2000_Sample/$exit
      -- CP-element group 154: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_length_2000_Sample/ack
      -- 
    ack_4019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_length_2148_2000_buf_ack_0, ack => outputPort_4_Daemon_CP_3687_elements(154)); -- 
    -- CP-element group 155:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	153 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (4) 
      -- CP-element group 155: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_length_2000_update_completed__ps
      -- CP-element group 155: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_length_2000_update_completed_
      -- CP-element group 155: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_length_2000_Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_active_packet_length_2000_Update/ack
      -- 
    ack_4024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_length_2148_2000_buf_ack_1, ack => outputPort_4_Daemon_CP_3687_elements(155)); -- 
    -- CP-element group 156:  join  transition  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	9 
    -- CP-element group 156: marked-predecessors 
    -- CP-element group 156: 	12 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	11 
    -- CP-element group 156:  members (1) 
      -- CP-element group 156: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_2001_sample_start_
      -- 
    outputPort_4_Daemon_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(9) & outputPort_4_Daemon_CP_3687_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  join  transition  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	9 
    -- CP-element group 157: marked-predecessors 
    -- CP-element group 157: 	176 
    -- CP-element group 157: 	179 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	14 
    -- CP-element group 157:  members (1) 
      -- CP-element group 157: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_2001_update_start_
      -- 
    outputPort_4_Daemon_cp_element_group_157: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_157"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(9) & outputPort_4_Daemon_CP_3687_elements(176) & outputPort_4_Daemon_CP_3687_elements(179);
      gj_outputPort_4_Daemon_cp_element_group_157 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(157), clk => clk, reset => reset); --
    end block;
    -- CP-element group 158:  join  transition  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	12 
    -- CP-element group 158:  members (1) 
      -- CP-element group 158: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_2001_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(158) is bound as output of CP function.
    -- CP-element group 159:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	14 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (1) 
      -- CP-element group 159: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_2001_update_start__ps
      -- 
    outputPort_4_Daemon_CP_3687_elements(159) <= outputPort_4_Daemon_CP_3687_elements(14);
    -- CP-element group 160:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	174 
    -- CP-element group 160: 	178 
    -- CP-element group 160: 	15 
    -- CP-element group 160:  members (2) 
      -- CP-element group 160: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_2001_update_completed__ps
      -- CP-element group 160: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_2001_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(160) is bound as output of CP function.
    -- CP-element group 161:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	7 
    -- CP-element group 161: successors 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_2001_loopback_trigger
      -- 
    outputPort_4_Daemon_CP_3687_elements(161) <= outputPort_4_Daemon_CP_3687_elements(7);
    -- CP-element group 162:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (2) 
      -- CP-element group 162: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_2001_loopback_sample_req_ps
      -- CP-element group 162: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_2001_loopback_sample_req
      -- 
    phi_stmt_2001_loopback_sample_req_4035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2001_loopback_sample_req_4035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(162), ack => phi_stmt_2001_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(162) is bound as output of CP function.
    -- CP-element group 163:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	8 
    -- CP-element group 163: successors 
    -- CP-element group 163:  members (1) 
      -- CP-element group 163: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_2001_entry_trigger
      -- 
    outputPort_4_Daemon_CP_3687_elements(163) <= outputPort_4_Daemon_CP_3687_elements(8);
    -- CP-element group 164:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (2) 
      -- CP-element group 164: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_2001_entry_sample_req
      -- CP-element group 164: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_2001_entry_sample_req_ps
      -- 
    phi_stmt_2001_entry_sample_req_4038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2001_entry_sample_req_4038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(164), ack => phi_stmt_2001_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(164) is bound as output of CP function.
    -- CP-element group 165:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: successors 
    -- CP-element group 165:  members (2) 
      -- CP-element group 165: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_2001_phi_mux_ack
      -- CP-element group 165: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/phi_stmt_2001_phi_mux_ack_ps
      -- 
    phi_stmt_2001_phi_mux_ack_4041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2001_ack_0, ack => outputPort_4_Daemon_CP_3687_elements(165)); -- 
    -- CP-element group 166:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: successors 
    -- CP-element group 166:  members (4) 
      -- CP-element group 166: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_2_2003_sample_start_
      -- CP-element group 166: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_2_2003_sample_completed_
      -- CP-element group 166: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_2_2003_sample_completed__ps
      -- CP-element group 166: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_2_2003_sample_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(166) is bound as output of CP function.
    -- CP-element group 167:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (2) 
      -- CP-element group 167: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_2_2003_update_start_
      -- CP-element group 167: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_2_2003_update_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(167) is bound as output of CP function.
    -- CP-element group 168:  join  transition  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	169 
    -- CP-element group 168: successors 
    -- CP-element group 168:  members (1) 
      -- CP-element group 168: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_2_2003_update_completed__ps
      -- 
    outputPort_4_Daemon_CP_3687_elements(168) <= outputPort_4_Daemon_CP_3687_elements(169);
    -- CP-element group 169:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	168 
    -- CP-element group 169:  members (1) 
      -- CP-element group 169: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_ZERO_2_2003_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(169) is a control-delay.
    cp_element_169_delay: control_delay_element  generic map(name => " 169_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_3687_elements(167), ack => outputPort_4_Daemon_CP_3687_elements(169), clk => clk, reset =>reset);
    -- CP-element group 170:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	172 
    -- CP-element group 170:  members (4) 
      -- CP-element group 170: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_priority_index_2004_sample_start__ps
      -- CP-element group 170: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_priority_index_2004_Sample/req
      -- CP-element group 170: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_priority_index_2004_Sample/$entry
      -- CP-element group 170: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_priority_index_2004_sample_start_
      -- 
    req_4062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(170), ack => next_priority_index_2103_2004_buf_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(170) is bound as output of CP function.
    -- CP-element group 171:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (4) 
      -- CP-element group 171: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_priority_index_2004_Update/req
      -- CP-element group 171: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_priority_index_2004_Update/$entry
      -- CP-element group 171: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_priority_index_2004_update_start_
      -- CP-element group 171: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_priority_index_2004_update_start__ps
      -- 
    req_4067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(171), ack => next_priority_index_2103_2004_buf_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(171) is bound as output of CP function.
    -- CP-element group 172:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	170 
    -- CP-element group 172: successors 
    -- CP-element group 172:  members (4) 
      -- CP-element group 172: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_priority_index_2004_Sample/ack
      -- CP-element group 172: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_priority_index_2004_sample_completed__ps
      -- CP-element group 172: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_priority_index_2004_Sample/$exit
      -- CP-element group 172: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_priority_index_2004_sample_completed_
      -- 
    ack_4063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_priority_index_2103_2004_buf_ack_0, ack => outputPort_4_Daemon_CP_3687_elements(172)); -- 
    -- CP-element group 173:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: successors 
    -- CP-element group 173:  members (4) 
      -- CP-element group 173: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_priority_index_2004_Update/ack
      -- CP-element group 173: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_priority_index_2004_Update/$exit
      -- CP-element group 173: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_priority_index_2004_update_completed_
      -- CP-element group 173: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/R_next_priority_index_2004_update_completed__ps
      -- 
    ack_4068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_priority_index_2103_2004_buf_ack_1, ack => outputPort_4_Daemon_CP_3687_elements(173)); -- 
    -- CP-element group 174:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	124 
    -- CP-element group 174: 	160 
    -- CP-element group 174: 	21 
    -- CP-element group 174: 	40 
    -- CP-element group 174: 	61 
    -- CP-element group 174: 	82 
    -- CP-element group 174: 	103 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	176 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/call_stmt_2032_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/call_stmt_2032_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/call_stmt_2032_Sample/crr
      -- 
    crr_4077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_4077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(174), ack => call_stmt_2032_call_req_0); -- 
    outputPort_4_Daemon_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(124) & outputPort_4_Daemon_CP_3687_elements(160) & outputPort_4_Daemon_CP_3687_elements(21) & outputPort_4_Daemon_CP_3687_elements(40) & outputPort_4_Daemon_CP_3687_elements(61) & outputPort_4_Daemon_CP_3687_elements(82) & outputPort_4_Daemon_CP_3687_elements(103);
      gj_outputPort_4_Daemon_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: marked-predecessors 
    -- CP-element group 175: 	177 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	177 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/call_stmt_2032_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/call_stmt_2032_update_start_
      -- CP-element group 175: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/call_stmt_2032_Update/ccr
      -- 
    ccr_4082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_4082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(175), ack => call_stmt_2032_call_req_1); -- 
    outputPort_4_Daemon_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= outputPort_4_Daemon_CP_3687_elements(177);
      gj_outputPort_4_Daemon_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	174 
    -- CP-element group 176: successors 
    -- CP-element group 176: marked-successors 
    -- CP-element group 176: 	157 
    -- CP-element group 176: 	120 
    -- CP-element group 176: 	17 
    -- CP-element group 176: 	36 
    -- CP-element group 176: 	57 
    -- CP-element group 176: 	78 
    -- CP-element group 176: 	99 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/call_stmt_2032_sample_completed_
      -- CP-element group 176: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/call_stmt_2032_Sample/cra
      -- CP-element group 176: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/call_stmt_2032_Sample/$exit
      -- 
    cra_4078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2032_call_ack_0, ack => outputPort_4_Daemon_CP_3687_elements(176)); -- 
    -- CP-element group 177:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	182 
    -- CP-element group 177: marked-successors 
    -- CP-element group 177: 	175 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/call_stmt_2032_Update/$exit
      -- CP-element group 177: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/call_stmt_2032_update_completed_
      -- CP-element group 177: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/call_stmt_2032_Update/cca
      -- 
    cca_4083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2032_call_ack_1, ack => outputPort_4_Daemon_CP_3687_elements(177)); -- 
    -- CP-element group 178:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	124 
    -- CP-element group 178: 	160 
    -- CP-element group 178: 	21 
    -- CP-element group 178: 	40 
    -- CP-element group 178: 	61 
    -- CP-element group 178: 	82 
    -- CP-element group 178: 	103 
    -- CP-element group 178: marked-predecessors 
    -- CP-element group 178: 	180 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/WPIPE_out_data_4_2257_Sample/req
      -- CP-element group 178: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/WPIPE_out_data_4_2257_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/WPIPE_out_data_4_2257_sample_start_
      -- 
    req_4091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(178), ack => WPIPE_out_data_4_2257_inst_req_0); -- 
    outputPort_4_Daemon_cp_element_group_178: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_178"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(124) & outputPort_4_Daemon_CP_3687_elements(160) & outputPort_4_Daemon_CP_3687_elements(21) & outputPort_4_Daemon_CP_3687_elements(40) & outputPort_4_Daemon_CP_3687_elements(61) & outputPort_4_Daemon_CP_3687_elements(82) & outputPort_4_Daemon_CP_3687_elements(103) & outputPort_4_Daemon_CP_3687_elements(180);
      gj_outputPort_4_Daemon_cp_element_group_178 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(178), clk => clk, reset => reset); --
    end block;
    -- CP-element group 179:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179: marked-successors 
    -- CP-element group 179: 	157 
    -- CP-element group 179: 	120 
    -- CP-element group 179: 	17 
    -- CP-element group 179: 	36 
    -- CP-element group 179: 	57 
    -- CP-element group 179: 	78 
    -- CP-element group 179: 	99 
    -- CP-element group 179:  members (6) 
      -- CP-element group 179: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/WPIPE_out_data_4_2257_Update/req
      -- CP-element group 179: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/WPIPE_out_data_4_2257_Update/$entry
      -- CP-element group 179: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/WPIPE_out_data_4_2257_Sample/ack
      -- CP-element group 179: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/WPIPE_out_data_4_2257_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/WPIPE_out_data_4_2257_update_start_
      -- CP-element group 179: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/WPIPE_out_data_4_2257_sample_completed_
      -- 
    ack_4092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_4_2257_inst_ack_0, ack => outputPort_4_Daemon_CP_3687_elements(179)); -- 
    req_4096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_3687_elements(179), ack => WPIPE_out_data_4_2257_inst_req_1); -- 
    -- CP-element group 180:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	182 
    -- CP-element group 180: marked-successors 
    -- CP-element group 180: 	178 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/WPIPE_out_data_4_2257_Update/ack
      -- CP-element group 180: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/WPIPE_out_data_4_2257_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/WPIPE_out_data_4_2257_update_completed_
      -- 
    ack_4097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_4_2257_inst_ack_1, ack => outputPort_4_Daemon_CP_3687_elements(180)); -- 
    -- CP-element group 181:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	9 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	10 
    -- CP-element group 181:  members (1) 
      -- CP-element group 181: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group outputPort_4_Daemon_CP_3687_elements(181) is a control-delay.
    cp_element_181_delay: control_delay_element  generic map(name => " 181_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_3687_elements(9), ack => outputPort_4_Daemon_CP_3687_elements(181), clk => clk, reset =>reset);
    -- CP-element group 182:  join  transition  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	177 
    -- CP-element group 182: 	180 
    -- CP-element group 182: 	12 
    -- CP-element group 182: 	13 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	6 
    -- CP-element group 182:  members (1) 
      -- CP-element group 182: 	 branch_block_stmt_1966/do_while_stmt_1967/do_while_stmt_1967_loop_body/$exit
      -- 
    outputPort_4_Daemon_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 7,2 => 7,3 => 7);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_3687_elements(177) & outputPort_4_Daemon_CP_3687_elements(180) & outputPort_4_Daemon_CP_3687_elements(12) & outputPort_4_Daemon_CP_3687_elements(13);
      gj_outputPort_4_Daemon_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  transition  input  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	5 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (2) 
      -- CP-element group 183: 	 branch_block_stmt_1966/do_while_stmt_1967/loop_exit/ack
      -- CP-element group 183: 	 branch_block_stmt_1966/do_while_stmt_1967/loop_exit/$exit
      -- 
    ack_4102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1967_branch_ack_0, ack => outputPort_4_Daemon_CP_3687_elements(183)); -- 
    -- CP-element group 184:  transition  input  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	5 
    -- CP-element group 184: successors 
    -- CP-element group 184:  members (2) 
      -- CP-element group 184: 	 branch_block_stmt_1966/do_while_stmt_1967/loop_taken/ack
      -- CP-element group 184: 	 branch_block_stmt_1966/do_while_stmt_1967/loop_taken/$exit
      -- 
    ack_4106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1967_branch_ack_1, ack => outputPort_4_Daemon_CP_3687_elements(184)); -- 
    -- CP-element group 185:  transition  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	3 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	1 
    -- CP-element group 185:  members (1) 
      -- CP-element group 185: 	 branch_block_stmt_1966/do_while_stmt_1967/$exit
      -- 
    outputPort_4_Daemon_CP_3687_elements(185) <= outputPort_4_Daemon_CP_3687_elements(3);
    outputPort_4_Daemon_do_while_stmt_1967_terminator_4107: loop_terminator -- 
      generic map (name => " outputPort_4_Daemon_do_while_stmt_1967_terminator_4107", max_iterations_in_flight =>7) 
      port map(loop_body_exit => outputPort_4_Daemon_CP_3687_elements(6),loop_continue => outputPort_4_Daemon_CP_3687_elements(184),loop_terminate => outputPort_4_Daemon_CP_3687_elements(183),loop_back => outputPort_4_Daemon_CP_3687_elements(4),loop_exit => outputPort_4_Daemon_CP_3687_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1969_phi_seq_3761_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_4_Daemon_CP_3687_elements(24);
      outputPort_4_Daemon_CP_3687_elements(27)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_4_Daemon_CP_3687_elements(27);
      outputPort_4_Daemon_CP_3687_elements(28)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_4_Daemon_CP_3687_elements(29);
      outputPort_4_Daemon_CP_3687_elements(25) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_4_Daemon_CP_3687_elements(22);
      outputPort_4_Daemon_CP_3687_elements(31)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_4_Daemon_CP_3687_elements(33);
      outputPort_4_Daemon_CP_3687_elements(32)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_4_Daemon_CP_3687_elements(34);
      outputPort_4_Daemon_CP_3687_elements(23) <= phi_mux_reqs(1);
      phi_stmt_1969_phi_seq_3761 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1969_phi_seq_3761") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_4_Daemon_CP_3687_elements(18), 
          phi_sample_ack => outputPort_4_Daemon_CP_3687_elements(19), 
          phi_update_req => outputPort_4_Daemon_CP_3687_elements(20), 
          phi_update_ack => outputPort_4_Daemon_CP_3687_elements(21), 
          phi_mux_ack => outputPort_4_Daemon_CP_3687_elements(26), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1973_phi_seq_3805_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_4_Daemon_CP_3687_elements(43);
      outputPort_4_Daemon_CP_3687_elements(46)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_4_Daemon_CP_3687_elements(46);
      outputPort_4_Daemon_CP_3687_elements(47)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_4_Daemon_CP_3687_elements(48);
      outputPort_4_Daemon_CP_3687_elements(44) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_4_Daemon_CP_3687_elements(41);
      outputPort_4_Daemon_CP_3687_elements(50)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_4_Daemon_CP_3687_elements(54);
      outputPort_4_Daemon_CP_3687_elements(51)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_4_Daemon_CP_3687_elements(55);
      outputPort_4_Daemon_CP_3687_elements(42) <= phi_mux_reqs(1);
      phi_stmt_1973_phi_seq_3805 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1973_phi_seq_3805") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_4_Daemon_CP_3687_elements(37), 
          phi_sample_ack => outputPort_4_Daemon_CP_3687_elements(38), 
          phi_update_req => outputPort_4_Daemon_CP_3687_elements(39), 
          phi_update_ack => outputPort_4_Daemon_CP_3687_elements(40), 
          phi_mux_ack => outputPort_4_Daemon_CP_3687_elements(45), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1978_phi_seq_3849_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_4_Daemon_CP_3687_elements(64);
      outputPort_4_Daemon_CP_3687_elements(67)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_4_Daemon_CP_3687_elements(67);
      outputPort_4_Daemon_CP_3687_elements(68)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_4_Daemon_CP_3687_elements(69);
      outputPort_4_Daemon_CP_3687_elements(65) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_4_Daemon_CP_3687_elements(62);
      outputPort_4_Daemon_CP_3687_elements(71)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_4_Daemon_CP_3687_elements(75);
      outputPort_4_Daemon_CP_3687_elements(72)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_4_Daemon_CP_3687_elements(76);
      outputPort_4_Daemon_CP_3687_elements(63) <= phi_mux_reqs(1);
      phi_stmt_1978_phi_seq_3849 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1978_phi_seq_3849") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_4_Daemon_CP_3687_elements(58), 
          phi_sample_ack => outputPort_4_Daemon_CP_3687_elements(59), 
          phi_update_req => outputPort_4_Daemon_CP_3687_elements(60), 
          phi_update_ack => outputPort_4_Daemon_CP_3687_elements(61), 
          phi_mux_ack => outputPort_4_Daemon_CP_3687_elements(66), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1983_phi_seq_3893_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_4_Daemon_CP_3687_elements(85);
      outputPort_4_Daemon_CP_3687_elements(88)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_4_Daemon_CP_3687_elements(88);
      outputPort_4_Daemon_CP_3687_elements(89)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_4_Daemon_CP_3687_elements(90);
      outputPort_4_Daemon_CP_3687_elements(86) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_4_Daemon_CP_3687_elements(83);
      outputPort_4_Daemon_CP_3687_elements(92)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_4_Daemon_CP_3687_elements(96);
      outputPort_4_Daemon_CP_3687_elements(93)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_4_Daemon_CP_3687_elements(97);
      outputPort_4_Daemon_CP_3687_elements(84) <= phi_mux_reqs(1);
      phi_stmt_1983_phi_seq_3893 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1983_phi_seq_3893") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_4_Daemon_CP_3687_elements(79), 
          phi_sample_ack => outputPort_4_Daemon_CP_3687_elements(80), 
          phi_update_req => outputPort_4_Daemon_CP_3687_elements(81), 
          phi_update_ack => outputPort_4_Daemon_CP_3687_elements(82), 
          phi_mux_ack => outputPort_4_Daemon_CP_3687_elements(87), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1988_phi_seq_3937_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_4_Daemon_CP_3687_elements(106);
      outputPort_4_Daemon_CP_3687_elements(109)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_4_Daemon_CP_3687_elements(109);
      outputPort_4_Daemon_CP_3687_elements(110)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_4_Daemon_CP_3687_elements(111);
      outputPort_4_Daemon_CP_3687_elements(107) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_4_Daemon_CP_3687_elements(104);
      outputPort_4_Daemon_CP_3687_elements(113)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_4_Daemon_CP_3687_elements(117);
      outputPort_4_Daemon_CP_3687_elements(114)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_4_Daemon_CP_3687_elements(118);
      outputPort_4_Daemon_CP_3687_elements(105) <= phi_mux_reqs(1);
      phi_stmt_1988_phi_seq_3937 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1988_phi_seq_3937") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_4_Daemon_CP_3687_elements(100), 
          phi_sample_ack => outputPort_4_Daemon_CP_3687_elements(101), 
          phi_update_req => outputPort_4_Daemon_CP_3687_elements(102), 
          phi_update_ack => outputPort_4_Daemon_CP_3687_elements(103), 
          phi_mux_ack => outputPort_4_Daemon_CP_3687_elements(108), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1993_phi_seq_3981_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_4_Daemon_CP_3687_elements(127);
      outputPort_4_Daemon_CP_3687_elements(130)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_4_Daemon_CP_3687_elements(130);
      outputPort_4_Daemon_CP_3687_elements(131)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_4_Daemon_CP_3687_elements(132);
      outputPort_4_Daemon_CP_3687_elements(128) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_4_Daemon_CP_3687_elements(125);
      outputPort_4_Daemon_CP_3687_elements(134)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_4_Daemon_CP_3687_elements(136);
      outputPort_4_Daemon_CP_3687_elements(135)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_4_Daemon_CP_3687_elements(137);
      outputPort_4_Daemon_CP_3687_elements(126) <= phi_mux_reqs(1);
      phi_stmt_1993_phi_seq_3981 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1993_phi_seq_3981") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_4_Daemon_CP_3687_elements(121), 
          phi_sample_ack => outputPort_4_Daemon_CP_3687_elements(122), 
          phi_update_req => outputPort_4_Daemon_CP_3687_elements(123), 
          phi_update_ack => outputPort_4_Daemon_CP_3687_elements(124), 
          phi_mux_ack => outputPort_4_Daemon_CP_3687_elements(129), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1997_phi_seq_4025_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_4_Daemon_CP_3687_elements(145);
      outputPort_4_Daemon_CP_3687_elements(148)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_4_Daemon_CP_3687_elements(148);
      outputPort_4_Daemon_CP_3687_elements(149)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_4_Daemon_CP_3687_elements(150);
      outputPort_4_Daemon_CP_3687_elements(146) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_4_Daemon_CP_3687_elements(143);
      outputPort_4_Daemon_CP_3687_elements(152)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_4_Daemon_CP_3687_elements(154);
      outputPort_4_Daemon_CP_3687_elements(153)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_4_Daemon_CP_3687_elements(155);
      outputPort_4_Daemon_CP_3687_elements(144) <= phi_mux_reqs(1);
      phi_stmt_1997_phi_seq_4025 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1997_phi_seq_4025") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_4_Daemon_CP_3687_elements(140), 
          phi_sample_ack => outputPort_4_Daemon_CP_3687_elements(141), 
          phi_update_req => outputPort_4_Daemon_CP_3687_elements(14), 
          phi_update_ack => outputPort_4_Daemon_CP_3687_elements(142), 
          phi_mux_ack => outputPort_4_Daemon_CP_3687_elements(147), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2001_phi_seq_4069_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_4_Daemon_CP_3687_elements(163);
      outputPort_4_Daemon_CP_3687_elements(166)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_4_Daemon_CP_3687_elements(166);
      outputPort_4_Daemon_CP_3687_elements(167)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_4_Daemon_CP_3687_elements(168);
      outputPort_4_Daemon_CP_3687_elements(164) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_4_Daemon_CP_3687_elements(161);
      outputPort_4_Daemon_CP_3687_elements(170)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_4_Daemon_CP_3687_elements(172);
      outputPort_4_Daemon_CP_3687_elements(171)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_4_Daemon_CP_3687_elements(173);
      outputPort_4_Daemon_CP_3687_elements(162) <= phi_mux_reqs(1);
      phi_stmt_2001_phi_seq_4069 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_2001_phi_seq_4069") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_4_Daemon_CP_3687_elements(11), 
          phi_sample_ack => outputPort_4_Daemon_CP_3687_elements(158), 
          phi_update_req => outputPort_4_Daemon_CP_3687_elements(159), 
          phi_update_ack => outputPort_4_Daemon_CP_3687_elements(160), 
          phi_mux_ack => outputPort_4_Daemon_CP_3687_elements(165), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3712_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= outputPort_4_Daemon_CP_3687_elements(7);
        preds(1)  <= outputPort_4_Daemon_CP_3687_elements(8);
        entry_tmerge_3712 : transition_merge -- 
          generic map(name => " entry_tmerge_3712")
          port map (preds => preds, symbol_out => outputPort_4_Daemon_CP_3687_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal EQ_u3_u1_2068_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2074_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2081_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2087_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2117_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2124_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2132_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2139_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2167_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2175_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2183_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2191_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2197_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2204_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2212_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2219_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2230_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2236_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2243_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2249_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_2110_wire : std_logic_vector(0 downto 0);
    signal MUX_2010_wire : std_logic_vector(7 downto 0);
    signal MUX_2014_wire : std_logic_vector(7 downto 0);
    signal MUX_2019_wire : std_logic_vector(7 downto 0);
    signal MUX_2023_wire : std_logic_vector(7 downto 0);
    signal MUX_2071_wire : std_logic_vector(0 downto 0);
    signal MUX_2077_wire : std_logic_vector(0 downto 0);
    signal MUX_2084_wire : std_logic_vector(0 downto 0);
    signal MUX_2090_wire : std_logic_vector(0 downto 0);
    signal MUX_2121_wire : std_logic_vector(7 downto 0);
    signal MUX_2128_wire : std_logic_vector(7 downto 0);
    signal MUX_2136_wire : std_logic_vector(7 downto 0);
    signal MUX_2143_wire : std_logic_vector(7 downto 0);
    signal MUX_2159_wire : std_logic_vector(7 downto 0);
    signal MUX_2201_wire : std_logic_vector(31 downto 0);
    signal MUX_2208_wire : std_logic_vector(31 downto 0);
    signal MUX_2216_wire : std_logic_vector(31 downto 0);
    signal MUX_2223_wire : std_logic_vector(31 downto 0);
    signal MUX_2233_wire : std_logic_vector(0 downto 0);
    signal MUX_2239_wire : std_logic_vector(0 downto 0);
    signal MUX_2246_wire : std_logic_vector(0 downto 0);
    signal MUX_2252_wire : std_logic_vector(0 downto 0);
    signal NEQ_u3_u1_2107_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_2164_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_2172_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_2180_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_2188_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_2078_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_2091_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_2240_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_2253_wire : std_logic_vector(0 downto 0);
    signal OR_u32_u32_2209_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_2224_wire : std_logic_vector(31 downto 0);
    signal OR_u8_u8_2015_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_2024_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_2129_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_2144_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_2145_wire : std_logic_vector(7 downto 0);
    signal RPIPE_noblock_obuf_1_4_1977_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_2_4_1982_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_3_4_1987_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_4_4_1992_wire : std_logic_vector(32 downto 0);
    signal R_ZERO_2_2003_wire_constant : std_logic_vector(1 downto 0);
    signal R_ZERO_33_1975_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1980_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1985_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1990_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_3_1995_wire_constant : std_logic_vector(2 downto 0);
    signal R_ZERO_8_1971_wire_constant : std_logic_vector(7 downto 0);
    signal R_ZERO_8_1999_wire_constant : std_logic_vector(7 downto 0);
    signal SUB_u8_u8_2153_wire : std_logic_vector(7 downto 0);
    signal SUB_u8_u8_2157_wire : std_logic_vector(7 downto 0);
    signal active_packet_1993 : std_logic_vector(2 downto 0);
    signal active_packet_length_1997 : std_logic_vector(7 downto 0);
    signal continue_2032 : std_logic_vector(0 downto 0);
    signal data_to_out_2226 : std_logic_vector(31 downto 0);
    signal down_counter_1969 : std_logic_vector(7 downto 0);
    signal konst_2008_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2009_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2012_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2013_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2017_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2018_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2021_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2022_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2028_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2035_wire_constant : std_logic_vector(32 downto 0);
    signal konst_2040_wire_constant : std_logic_vector(32 downto 0);
    signal konst_2045_wire_constant : std_logic_vector(32 downto 0);
    signal konst_2050_wire_constant : std_logic_vector(32 downto 0);
    signal konst_2067_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2070_wire_constant : std_logic_vector(0 downto 0);
    signal konst_2073_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2076_wire_constant : std_logic_vector(0 downto 0);
    signal konst_2080_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2083_wire_constant : std_logic_vector(0 downto 0);
    signal konst_2086_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2089_wire_constant : std_logic_vector(0 downto 0);
    signal konst_2106_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2109_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2116_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2120_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2123_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2127_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2131_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2135_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2138_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2142_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2152_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2156_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2166_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2174_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2182_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2190_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2196_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2200_wire_constant : std_logic_vector(31 downto 0);
    signal konst_2203_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2207_wire_constant : std_logic_vector(31 downto 0);
    signal konst_2211_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2215_wire_constant : std_logic_vector(31 downto 0);
    signal konst_2218_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2222_wire_constant : std_logic_vector(31 downto 0);
    signal konst_2229_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2232_wire_constant : std_logic_vector(0 downto 0);
    signal konst_2235_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2238_wire_constant : std_logic_vector(0 downto 0);
    signal konst_2242_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2245_wire_constant : std_logic_vector(0 downto 0);
    signal konst_2248_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2251_wire_constant : std_logic_vector(0 downto 0);
    signal konst_2270_wire_constant : std_logic_vector(0 downto 0);
    signal next_active_packet_2103 : std_logic_vector(2 downto 0);
    signal next_active_packet_2103_1996_buffered : std_logic_vector(2 downto 0);
    signal next_active_packet_length_2148 : std_logic_vector(7 downto 0);
    signal next_active_packet_length_2148_2000_buffered : std_logic_vector(7 downto 0);
    signal next_down_counter_2161 : std_logic_vector(7 downto 0);
    signal next_down_counter_2161_1972_buffered : std_logic_vector(7 downto 0);
    signal next_priority_index_2103 : std_logic_vector(1 downto 0);
    signal next_priority_index_2103_2004_buffered : std_logic_vector(1 downto 0);
    signal p1_valid_2037 : std_logic_vector(0 downto 0);
    signal p2_valid_2042 : std_logic_vector(0 downto 0);
    signal p3_valid_2047 : std_logic_vector(0 downto 0);
    signal p4_valid_2052 : std_logic_vector(0 downto 0);
    signal pkt_1_e_word_1973 : std_logic_vector(32 downto 0);
    signal pkt_2_e_word_1978 : std_logic_vector(32 downto 0);
    signal pkt_3_e_word_1983 : std_logic_vector(32 downto 0);
    signal pkt_4_e_word_1988 : std_logic_vector(32 downto 0);
    signal priority_index_2001 : std_logic_vector(1 downto 0);
    signal read_from_1_2169 : std_logic_vector(0 downto 0);
    signal read_from_2_2177 : std_logic_vector(0 downto 0);
    signal read_from_3_2185 : std_logic_vector(0 downto 0);
    signal read_from_4_2193 : std_logic_vector(0 downto 0);
    signal send_flag_2255 : std_logic_vector(0 downto 0);
    signal senderPort_2026 : std_logic_vector(7 downto 0);
    signal slice_2119_wire : std_logic_vector(7 downto 0);
    signal slice_2126_wire : std_logic_vector(7 downto 0);
    signal slice_2134_wire : std_logic_vector(7 downto 0);
    signal slice_2141_wire : std_logic_vector(7 downto 0);
    signal slice_2199_wire : std_logic_vector(31 downto 0);
    signal slice_2206_wire : std_logic_vector(31 downto 0);
    signal slice_2214_wire : std_logic_vector(31 downto 0);
    signal slice_2221_wire : std_logic_vector(31 downto 0);
    signal started_new_packet_2112 : std_logic_vector(0 downto 0);
    signal type_cast_2030_wire_constant : std_logic_vector(0 downto 0);
    signal valid_active_pkt_word_read_2093 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_ZERO_2_2003_wire_constant <= "00";
    R_ZERO_33_1975_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1980_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1985_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1990_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_3_1995_wire_constant <= "000";
    R_ZERO_8_1971_wire_constant <= "00000000";
    R_ZERO_8_1999_wire_constant <= "00000000";
    konst_2008_wire_constant <= "00000000";
    konst_2009_wire_constant <= "00000000";
    konst_2012_wire_constant <= "00000001";
    konst_2013_wire_constant <= "00000000";
    konst_2017_wire_constant <= "00000010";
    konst_2018_wire_constant <= "00000000";
    konst_2021_wire_constant <= "00000011";
    konst_2022_wire_constant <= "00000000";
    konst_2028_wire_constant <= "00000011";
    konst_2035_wire_constant <= "000000000000000000000000000100000";
    konst_2040_wire_constant <= "000000000000000000000000000100000";
    konst_2045_wire_constant <= "000000000000000000000000000100000";
    konst_2050_wire_constant <= "000000000000000000000000000100000";
    konst_2067_wire_constant <= "001";
    konst_2070_wire_constant <= "0";
    konst_2073_wire_constant <= "010";
    konst_2076_wire_constant <= "0";
    konst_2080_wire_constant <= "011";
    konst_2083_wire_constant <= "0";
    konst_2086_wire_constant <= "100";
    konst_2089_wire_constant <= "0";
    konst_2106_wire_constant <= "000";
    konst_2109_wire_constant <= "00000000";
    konst_2116_wire_constant <= "001";
    konst_2120_wire_constant <= "00000000";
    konst_2123_wire_constant <= "010";
    konst_2127_wire_constant <= "00000000";
    konst_2131_wire_constant <= "011";
    konst_2135_wire_constant <= "00000000";
    konst_2138_wire_constant <= "100";
    konst_2142_wire_constant <= "00000000";
    konst_2152_wire_constant <= "00000001";
    konst_2156_wire_constant <= "00000001";
    konst_2166_wire_constant <= "001";
    konst_2174_wire_constant <= "010";
    konst_2182_wire_constant <= "011";
    konst_2190_wire_constant <= "100";
    konst_2196_wire_constant <= "001";
    konst_2200_wire_constant <= "00000000000000000000000000000000";
    konst_2203_wire_constant <= "010";
    konst_2207_wire_constant <= "00000000000000000000000000000000";
    konst_2211_wire_constant <= "011";
    konst_2215_wire_constant <= "00000000000000000000000000000000";
    konst_2218_wire_constant <= "100";
    konst_2222_wire_constant <= "00000000000000000000000000000000";
    konst_2229_wire_constant <= "001";
    konst_2232_wire_constant <= "0";
    konst_2235_wire_constant <= "010";
    konst_2238_wire_constant <= "0";
    konst_2242_wire_constant <= "011";
    konst_2245_wire_constant <= "0";
    konst_2248_wire_constant <= "100";
    konst_2251_wire_constant <= "0";
    konst_2270_wire_constant <= "1";
    type_cast_2030_wire_constant <= "0";
    phi_stmt_1969: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_8_1971_wire_constant & next_down_counter_2161_1972_buffered;
      req <= phi_stmt_1969_req_0 & phi_stmt_1969_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1969",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1969_ack_0,
          idata => idata,
          odata => down_counter_1969,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1969
    phi_stmt_1973: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1975_wire_constant & RPIPE_noblock_obuf_1_4_1977_wire;
      req <= phi_stmt_1973_req_0 & phi_stmt_1973_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1973",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1973_ack_0,
          idata => idata,
          odata => pkt_1_e_word_1973,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1973
    phi_stmt_1978: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1980_wire_constant & RPIPE_noblock_obuf_2_4_1982_wire;
      req <= phi_stmt_1978_req_0 & phi_stmt_1978_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1978",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1978_ack_0,
          idata => idata,
          odata => pkt_2_e_word_1978,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1978
    phi_stmt_1983: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1985_wire_constant & RPIPE_noblock_obuf_3_4_1987_wire;
      req <= phi_stmt_1983_req_0 & phi_stmt_1983_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1983",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1983_ack_0,
          idata => idata,
          odata => pkt_3_e_word_1983,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1983
    phi_stmt_1988: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1990_wire_constant & RPIPE_noblock_obuf_4_4_1992_wire;
      req <= phi_stmt_1988_req_0 & phi_stmt_1988_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1988",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1988_ack_0,
          idata => idata,
          odata => pkt_4_e_word_1988,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1988
    phi_stmt_1993: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_3_1995_wire_constant & next_active_packet_2103_1996_buffered;
      req <= phi_stmt_1993_req_0 & phi_stmt_1993_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1993",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1993_ack_0,
          idata => idata,
          odata => active_packet_1993,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1993
    phi_stmt_1997: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_8_1999_wire_constant & next_active_packet_length_2148_2000_buffered;
      req <= phi_stmt_1997_req_0 & phi_stmt_1997_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1997",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1997_ack_0,
          idata => idata,
          odata => active_packet_length_1997,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1997
    phi_stmt_2001: Block -- phi operator 
      signal idata: std_logic_vector(3 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_2_2003_wire_constant & next_priority_index_2103_2004_buffered;
      req <= phi_stmt_2001_req_0 & phi_stmt_2001_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2001",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 2) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2001_ack_0,
          idata => idata,
          odata => priority_index_2001,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2001
    -- flow-through select operator MUX_2010_inst
    MUX_2010_wire <= konst_2008_wire_constant when (read_from_1_2169(0) /=  '0') else konst_2009_wire_constant;
    -- flow-through select operator MUX_2014_inst
    MUX_2014_wire <= konst_2012_wire_constant when (read_from_2_2177(0) /=  '0') else konst_2013_wire_constant;
    -- flow-through select operator MUX_2019_inst
    MUX_2019_wire <= konst_2017_wire_constant when (read_from_3_2185(0) /=  '0') else konst_2018_wire_constant;
    -- flow-through select operator MUX_2023_inst
    MUX_2023_wire <= konst_2021_wire_constant when (read_from_4_2193(0) /=  '0') else konst_2022_wire_constant;
    -- flow-through select operator MUX_2071_inst
    MUX_2071_wire <= p1_valid_2037 when (EQ_u3_u1_2068_wire(0) /=  '0') else konst_2070_wire_constant;
    -- flow-through select operator MUX_2077_inst
    MUX_2077_wire <= p2_valid_2042 when (EQ_u3_u1_2074_wire(0) /=  '0') else konst_2076_wire_constant;
    -- flow-through select operator MUX_2084_inst
    MUX_2084_wire <= p3_valid_2047 when (EQ_u3_u1_2081_wire(0) /=  '0') else konst_2083_wire_constant;
    -- flow-through select operator MUX_2090_inst
    MUX_2090_wire <= p4_valid_2052 when (EQ_u3_u1_2087_wire(0) /=  '0') else konst_2089_wire_constant;
    -- flow-through select operator MUX_2121_inst
    MUX_2121_wire <= slice_2119_wire when (EQ_u3_u1_2117_wire(0) /=  '0') else konst_2120_wire_constant;
    -- flow-through select operator MUX_2128_inst
    MUX_2128_wire <= slice_2126_wire when (EQ_u3_u1_2124_wire(0) /=  '0') else konst_2127_wire_constant;
    -- flow-through select operator MUX_2136_inst
    MUX_2136_wire <= slice_2134_wire when (EQ_u3_u1_2132_wire(0) /=  '0') else konst_2135_wire_constant;
    -- flow-through select operator MUX_2143_inst
    MUX_2143_wire <= slice_2141_wire when (EQ_u3_u1_2139_wire(0) /=  '0') else konst_2142_wire_constant;
    -- flow-through select operator MUX_2147_inst
    next_active_packet_length_2148 <= OR_u8_u8_2145_wire when (started_new_packet_2112(0) /=  '0') else active_packet_length_1997;
    -- flow-through select operator MUX_2159_inst
    MUX_2159_wire <= SUB_u8_u8_2157_wire when (valid_active_pkt_word_read_2093(0) /=  '0') else down_counter_1969;
    -- flow-through select operator MUX_2160_inst
    next_down_counter_2161 <= SUB_u8_u8_2153_wire when (started_new_packet_2112(0) /=  '0') else MUX_2159_wire;
    -- flow-through select operator MUX_2201_inst
    MUX_2201_wire <= slice_2199_wire when (EQ_u3_u1_2197_wire(0) /=  '0') else konst_2200_wire_constant;
    -- flow-through select operator MUX_2208_inst
    MUX_2208_wire <= slice_2206_wire when (EQ_u3_u1_2204_wire(0) /=  '0') else konst_2207_wire_constant;
    -- flow-through select operator MUX_2216_inst
    MUX_2216_wire <= slice_2214_wire when (EQ_u3_u1_2212_wire(0) /=  '0') else konst_2215_wire_constant;
    -- flow-through select operator MUX_2223_inst
    MUX_2223_wire <= slice_2221_wire when (EQ_u3_u1_2219_wire(0) /=  '0') else konst_2222_wire_constant;
    -- flow-through select operator MUX_2233_inst
    MUX_2233_wire <= p1_valid_2037 when (EQ_u3_u1_2230_wire(0) /=  '0') else konst_2232_wire_constant;
    -- flow-through select operator MUX_2239_inst
    MUX_2239_wire <= p2_valid_2042 when (EQ_u3_u1_2236_wire(0) /=  '0') else konst_2238_wire_constant;
    -- flow-through select operator MUX_2246_inst
    MUX_2246_wire <= p3_valid_2047 when (EQ_u3_u1_2243_wire(0) /=  '0') else konst_2245_wire_constant;
    -- flow-through select operator MUX_2252_inst
    MUX_2252_wire <= p4_valid_2052 when (EQ_u3_u1_2249_wire(0) /=  '0') else konst_2251_wire_constant;
    -- flow-through slice operator slice_2119_inst
    slice_2119_wire <= pkt_1_e_word_1973(15 downto 8);
    -- flow-through slice operator slice_2126_inst
    slice_2126_wire <= pkt_2_e_word_1978(15 downto 8);
    -- flow-through slice operator slice_2134_inst
    slice_2134_wire <= pkt_3_e_word_1983(15 downto 8);
    -- flow-through slice operator slice_2141_inst
    slice_2141_wire <= pkt_4_e_word_1988(15 downto 8);
    -- flow-through slice operator slice_2199_inst
    slice_2199_wire <= pkt_1_e_word_1973(31 downto 0);
    -- flow-through slice operator slice_2206_inst
    slice_2206_wire <= pkt_2_e_word_1978(31 downto 0);
    -- flow-through slice operator slice_2214_inst
    slice_2214_wire <= pkt_3_e_word_1983(31 downto 0);
    -- flow-through slice operator slice_2221_inst
    slice_2221_wire <= pkt_4_e_word_1988(31 downto 0);
    next_active_packet_2103_1996_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_active_packet_2103_1996_buf_req_0;
      next_active_packet_2103_1996_buf_ack_0<= wack(0);
      rreq(0) <= next_active_packet_2103_1996_buf_req_1;
      next_active_packet_2103_1996_buf_ack_1<= rack(0);
      next_active_packet_2103_1996_buf : InterlockBuffer generic map ( -- 
        name => "next_active_packet_2103_1996_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_active_packet_2103,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_active_packet_2103_1996_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_active_packet_length_2148_2000_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_active_packet_length_2148_2000_buf_req_0;
      next_active_packet_length_2148_2000_buf_ack_0<= wack(0);
      rreq(0) <= next_active_packet_length_2148_2000_buf_req_1;
      next_active_packet_length_2148_2000_buf_ack_1<= rack(0);
      next_active_packet_length_2148_2000_buf : InterlockBuffer generic map ( -- 
        name => "next_active_packet_length_2148_2000_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_active_packet_length_2148,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_active_packet_length_2148_2000_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_down_counter_2161_1972_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_down_counter_2161_1972_buf_req_0;
      next_down_counter_2161_1972_buf_ack_0<= wack(0);
      rreq(0) <= next_down_counter_2161_1972_buf_req_1;
      next_down_counter_2161_1972_buf_ack_1<= rack(0);
      next_down_counter_2161_1972_buf : InterlockBuffer generic map ( -- 
        name => "next_down_counter_2161_1972_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_down_counter_2161,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_down_counter_2161_1972_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_priority_index_2103_2004_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_priority_index_2103_2004_buf_req_0;
      next_priority_index_2103_2004_buf_ack_0<= wack(0);
      rreq(0) <= next_priority_index_2103_2004_buf_req_1;
      next_priority_index_2103_2004_buf_ack_1<= rack(0);
      next_priority_index_2103_2004_buf : InterlockBuffer generic map ( -- 
        name => "next_priority_index_2103_2004_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 2,
        out_data_width => 2,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_priority_index_2103,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_priority_index_2103_2004_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1967_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_2270_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1967_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1967_branch_req_0,
          ack0 => do_while_stmt_1967_branch_ack_0,
          ack1 => do_while_stmt_1967_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- flow through binary operator AND_u1_u1_2111_inst
    started_new_packet_2112 <= (NEQ_u3_u1_2107_wire and EQ_u8_u1_2110_wire);
    -- flow through binary operator BITSEL_u33_u1_2036_inst
    process(pkt_1_e_word_1973) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_1_e_word_1973, konst_2035_wire_constant, tmp_var);
      p1_valid_2037 <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u33_u1_2041_inst
    process(pkt_2_e_word_1978) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_2_e_word_1978, konst_2040_wire_constant, tmp_var);
      p2_valid_2042 <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u33_u1_2046_inst
    process(pkt_3_e_word_1983) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_3_e_word_1983, konst_2045_wire_constant, tmp_var);
      p3_valid_2047 <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u33_u1_2051_inst
    process(pkt_4_e_word_1988) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_4_e_word_1988, konst_2050_wire_constant, tmp_var);
      p4_valid_2052 <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_2068_inst
    process(active_packet_1993) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1993, konst_2067_wire_constant, tmp_var);
      EQ_u3_u1_2068_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_2074_inst
    process(active_packet_1993) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1993, konst_2073_wire_constant, tmp_var);
      EQ_u3_u1_2074_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_2081_inst
    process(active_packet_1993) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1993, konst_2080_wire_constant, tmp_var);
      EQ_u3_u1_2081_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_2087_inst
    process(active_packet_1993) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1993, konst_2086_wire_constant, tmp_var);
      EQ_u3_u1_2087_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_2117_inst
    process(next_active_packet_2103) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_2103, konst_2116_wire_constant, tmp_var);
      EQ_u3_u1_2117_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_2124_inst
    process(next_active_packet_2103) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_2103, konst_2123_wire_constant, tmp_var);
      EQ_u3_u1_2124_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_2132_inst
    process(next_active_packet_2103) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_2103, konst_2131_wire_constant, tmp_var);
      EQ_u3_u1_2132_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_2139_inst
    process(next_active_packet_2103) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_2103, konst_2138_wire_constant, tmp_var);
      EQ_u3_u1_2139_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_2167_inst
    process(next_active_packet_2103) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_2103, konst_2166_wire_constant, tmp_var);
      EQ_u3_u1_2167_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_2175_inst
    process(next_active_packet_2103) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_2103, konst_2174_wire_constant, tmp_var);
      EQ_u3_u1_2175_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_2183_inst
    process(next_active_packet_2103) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_2103, konst_2182_wire_constant, tmp_var);
      EQ_u3_u1_2183_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_2191_inst
    process(next_active_packet_2103) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_2103, konst_2190_wire_constant, tmp_var);
      EQ_u3_u1_2191_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_2197_inst
    process(next_active_packet_2103) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_2103, konst_2196_wire_constant, tmp_var);
      EQ_u3_u1_2197_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_2204_inst
    process(next_active_packet_2103) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_2103, konst_2203_wire_constant, tmp_var);
      EQ_u3_u1_2204_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_2212_inst
    process(next_active_packet_2103) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_2103, konst_2211_wire_constant, tmp_var);
      EQ_u3_u1_2212_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_2219_inst
    process(next_active_packet_2103) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_2103, konst_2218_wire_constant, tmp_var);
      EQ_u3_u1_2219_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_2230_inst
    process(next_active_packet_2103) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_2103, konst_2229_wire_constant, tmp_var);
      EQ_u3_u1_2230_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_2236_inst
    process(next_active_packet_2103) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_2103, konst_2235_wire_constant, tmp_var);
      EQ_u3_u1_2236_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_2243_inst
    process(next_active_packet_2103) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_2103, konst_2242_wire_constant, tmp_var);
      EQ_u3_u1_2243_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_2249_inst
    process(next_active_packet_2103) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_2103, konst_2248_wire_constant, tmp_var);
      EQ_u3_u1_2249_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u8_u1_2110_inst
    process(down_counter_1969) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(down_counter_1969, konst_2109_wire_constant, tmp_var);
      EQ_u8_u1_2110_wire <= tmp_var; --
    end process;
    -- flow through binary operator NEQ_u3_u1_2107_inst
    process(next_active_packet_2103) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(next_active_packet_2103, konst_2106_wire_constant, tmp_var);
      NEQ_u3_u1_2107_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_2164_inst
    process(p1_valid_2037) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p1_valid_2037, tmp_var);
      NOT_u1_u1_2164_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_2172_inst
    process(p2_valid_2042) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p2_valid_2042, tmp_var);
      NOT_u1_u1_2172_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_2180_inst
    process(p3_valid_2047) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p3_valid_2047, tmp_var);
      NOT_u1_u1_2180_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_2188_inst
    process(p4_valid_2052) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p4_valid_2052, tmp_var);
      NOT_u1_u1_2188_wire <= tmp_var; -- 
    end process;
    -- flow through binary operator OR_u1_u1_2078_inst
    OR_u1_u1_2078_wire <= (MUX_2071_wire or MUX_2077_wire);
    -- flow through binary operator OR_u1_u1_2091_inst
    OR_u1_u1_2091_wire <= (MUX_2084_wire or MUX_2090_wire);
    -- flow through binary operator OR_u1_u1_2092_inst
    valid_active_pkt_word_read_2093 <= (OR_u1_u1_2078_wire or OR_u1_u1_2091_wire);
    -- flow through binary operator OR_u1_u1_2168_inst
    read_from_1_2169 <= (NOT_u1_u1_2164_wire or EQ_u3_u1_2167_wire);
    -- flow through binary operator OR_u1_u1_2176_inst
    read_from_2_2177 <= (NOT_u1_u1_2172_wire or EQ_u3_u1_2175_wire);
    -- flow through binary operator OR_u1_u1_2184_inst
    read_from_3_2185 <= (NOT_u1_u1_2180_wire or EQ_u3_u1_2183_wire);
    -- flow through binary operator OR_u1_u1_2192_inst
    read_from_4_2193 <= (NOT_u1_u1_2188_wire or EQ_u3_u1_2191_wire);
    -- flow through binary operator OR_u1_u1_2240_inst
    OR_u1_u1_2240_wire <= (MUX_2233_wire or MUX_2239_wire);
    -- flow through binary operator OR_u1_u1_2253_inst
    OR_u1_u1_2253_wire <= (MUX_2246_wire or MUX_2252_wire);
    -- flow through binary operator OR_u1_u1_2254_inst
    send_flag_2255 <= (OR_u1_u1_2240_wire or OR_u1_u1_2253_wire);
    -- flow through binary operator OR_u32_u32_2209_inst
    OR_u32_u32_2209_wire <= (MUX_2201_wire or MUX_2208_wire);
    -- flow through binary operator OR_u32_u32_2224_inst
    OR_u32_u32_2224_wire <= (MUX_2216_wire or MUX_2223_wire);
    -- flow through binary operator OR_u32_u32_2225_inst
    data_to_out_2226 <= (OR_u32_u32_2209_wire or OR_u32_u32_2224_wire);
    -- flow through binary operator OR_u8_u8_2015_inst
    OR_u8_u8_2015_wire <= (MUX_2010_wire or MUX_2014_wire);
    -- flow through binary operator OR_u8_u8_2024_inst
    OR_u8_u8_2024_wire <= (MUX_2019_wire or MUX_2023_wire);
    -- flow through binary operator OR_u8_u8_2025_inst
    senderPort_2026 <= (OR_u8_u8_2015_wire or OR_u8_u8_2024_wire);
    -- flow through binary operator OR_u8_u8_2129_inst
    OR_u8_u8_2129_wire <= (MUX_2121_wire or MUX_2128_wire);
    -- flow through binary operator OR_u8_u8_2144_inst
    OR_u8_u8_2144_wire <= (MUX_2136_wire or MUX_2143_wire);
    -- flow through binary operator OR_u8_u8_2145_inst
    OR_u8_u8_2145_wire <= (OR_u8_u8_2129_wire or OR_u8_u8_2144_wire);
    -- flow through binary operator SUB_u8_u8_2153_inst
    SUB_u8_u8_2153_wire <= std_logic_vector(unsigned(next_active_packet_length_2148) - unsigned(konst_2152_wire_constant));
    -- flow through binary operator SUB_u8_u8_2157_inst
    SUB_u8_u8_2157_wire <= std_logic_vector(unsigned(down_counter_1969) - unsigned(konst_2156_wire_constant));
    -- shared inport operator group (0) : RPIPE_noblock_obuf_1_4_1977_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_1_4_1977_inst_req_0;
      RPIPE_noblock_obuf_1_4_1977_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_1_4_1977_inst_req_1;
      RPIPE_noblock_obuf_1_4_1977_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_1_2169(0);
      RPIPE_noblock_obuf_1_4_1977_wire <= data_out(32 downto 0);
      noblock_obuf_1_4_read_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_4_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_4_read_0: InputPortRevised -- 
        generic map ( name => "noblock_obuf_1_4_read_0", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_1_4_pipe_read_req(0),
          oack => noblock_obuf_1_4_pipe_read_ack(0),
          odata => noblock_obuf_1_4_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_noblock_obuf_2_4_1982_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_2_4_1982_inst_req_0;
      RPIPE_noblock_obuf_2_4_1982_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_2_4_1982_inst_req_1;
      RPIPE_noblock_obuf_2_4_1982_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_2_2177(0);
      RPIPE_noblock_obuf_2_4_1982_wire <= data_out(32 downto 0);
      noblock_obuf_2_4_read_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_4_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_4_read_1: InputPortRevised -- 
        generic map ( name => "noblock_obuf_2_4_read_1", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_2_4_pipe_read_req(0),
          oack => noblock_obuf_2_4_pipe_read_ack(0),
          odata => noblock_obuf_2_4_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_noblock_obuf_3_4_1987_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_3_4_1987_inst_req_0;
      RPIPE_noblock_obuf_3_4_1987_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_3_4_1987_inst_req_1;
      RPIPE_noblock_obuf_3_4_1987_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_3_2185(0);
      RPIPE_noblock_obuf_3_4_1987_wire <= data_out(32 downto 0);
      noblock_obuf_3_4_read_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_4_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_4_read_2: InputPortRevised -- 
        generic map ( name => "noblock_obuf_3_4_read_2", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_3_4_pipe_read_req(0),
          oack => noblock_obuf_3_4_pipe_read_ack(0),
          odata => noblock_obuf_3_4_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_noblock_obuf_4_4_1992_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_4_4_1992_inst_req_0;
      RPIPE_noblock_obuf_4_4_1992_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_4_4_1992_inst_req_1;
      RPIPE_noblock_obuf_4_4_1992_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_4_2193(0);
      RPIPE_noblock_obuf_4_4_1992_wire <= data_out(32 downto 0);
      noblock_obuf_4_4_read_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_4_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_4_read_3: InputPortRevised -- 
        generic map ( name => "noblock_obuf_4_4_read_3", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_4_4_pipe_read_req(0),
          oack => noblock_obuf_4_4_pipe_read_ack(0),
          odata => noblock_obuf_4_4_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_out_data_4_2257_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_out_data_4_2257_inst_req_0;
      WPIPE_out_data_4_2257_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_out_data_4_2257_inst_req_1;
      WPIPE_out_data_4_2257_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_flag_2255(0);
      data_in <= data_to_out_2226;
      out_data_4_write_0_gI: SplitGuardInterface generic map(name => "out_data_4_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      out_data_4_write_0: OutputPortRevised -- 
        generic map ( name => "out_data_4", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => out_data_4_pipe_write_req(0),
          oack => out_data_4_pipe_write_ack(0),
          odata => out_data_4_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_2032_call 
    updateCounter_call_group_0: Block -- 
      signal data_in: std_logic_vector(16 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2032_call_req_0;
      call_stmt_2032_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2032_call_req_1;
      call_stmt_2032_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      updateCounter_call_group_0_gI: SplitGuardInterface generic map(name => "updateCounter_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= senderPort_2026 & konst_2028_wire_constant & type_cast_2030_wire_constant;
      continue_2032 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 17,
        owidth => 17,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => updateCounter_call_reqs(0),
          ackR => updateCounter_call_acks(0),
          dataR => updateCounter_call_data(16 downto 0),
          tagR => updateCounter_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => updateCounter_return_acks(0), -- cross-over
          ackL => updateCounter_return_reqs(0), -- cross-over
          dataL => updateCounter_return_data(0 downto 0),
          tagL => updateCounter_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    volatile_operator_prioritySelect_6468: prioritySelect_Volatile port map(down_counter => down_counter_1969, active_packet => active_packet_1993, priority_index => priority_index_2001, p1_valid => p1_valid_2037, p2_valid => p2_valid_2042, p3_valid => p3_valid_2047, p4_valid => p4_valid_2052, next_active_packet => next_active_packet_2103, next_priority_index => next_priority_index_2103); 
    -- 
  end Block; -- data_path
  -- 
end outputPort_4_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity prioritySelect_Volatile is -- 
  port ( -- 
    down_counter : in  std_logic_vector(7 downto 0);
    active_packet : in  std_logic_vector(2 downto 0);
    priority_index : in  std_logic_vector(1 downto 0);
    p1_valid : in  std_logic_vector(0 downto 0);
    p2_valid : in  std_logic_vector(0 downto 0);
    p3_valid : in  std_logic_vector(0 downto 0);
    p4_valid : in  std_logic_vector(0 downto 0);
    next_active_packet : out  std_logic_vector(2 downto 0);
    next_priority_index : out  std_logic_vector(1 downto 0)-- 
  );
  -- 
end entity prioritySelect_Volatile;
architecture prioritySelect_Volatile_arch of prioritySelect_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(17-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal down_counter_buffer :  std_logic_vector(7 downto 0);
  signal active_packet_buffer :  std_logic_vector(2 downto 0);
  signal priority_index_buffer :  std_logic_vector(1 downto 0);
  signal p1_valid_buffer :  std_logic_vector(0 downto 0);
  signal p2_valid_buffer :  std_logic_vector(0 downto 0);
  signal p3_valid_buffer :  std_logic_vector(0 downto 0);
  signal p4_valid_buffer :  std_logic_vector(0 downto 0);
  -- output port buffer signals
  signal next_active_packet_buffer :  std_logic_vector(2 downto 0);
  signal next_priority_index_buffer :  std_logic_vector(1 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  down_counter_buffer <= down_counter;
  active_packet_buffer <= active_packet;
  priority_index_buffer <= priority_index;
  p1_valid_buffer <= p1_valid;
  p2_valid_buffer <= p2_valid;
  p3_valid_buffer <= p3_valid;
  p4_valid_buffer <= p4_valid;
  -- output handling  -------------------------------------------------------
  next_active_packet <= next_active_packet_buffer;
  next_priority_index <= next_priority_index_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal ADD_u2_u2_1002_wire : std_logic_vector(1 downto 0);
    signal ADD_u2_u2_1020_wire : std_logic_vector(1 downto 0);
    signal ADD_u2_u2_1024_wire : std_logic_vector(1 downto 0);
    signal ADD_u2_u2_1028_wire : std_logic_vector(1 downto 0);
    signal ADD_u2_u2_1032_wire : std_logic_vector(1 downto 0);
    signal ADD_u2_u2_986_wire : std_logic_vector(1 downto 0);
    signal ADD_u2_u2_994_wire : std_logic_vector(1 downto 0);
    signal ADD_u3_u3_1005_wire : std_logic_vector(2 downto 0);
    signal ADD_u3_u3_981_wire : std_logic_vector(2 downto 0);
    signal ADD_u3_u3_989_wire : std_logic_vector(2 downto 0);
    signal ADD_u3_u3_997_wire : std_logic_vector(2 downto 0);
    signal CONCAT_u1_u3_1003_wire : std_logic_vector(2 downto 0);
    signal CONCAT_u1_u3_979_wire : std_logic_vector(2 downto 0);
    signal CONCAT_u1_u3_987_wire : std_logic_vector(2 downto 0);
    signal CONCAT_u1_u3_995_wire : std_logic_vector(2 downto 0);
    signal EQ_u2_u1_839_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_845_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_852_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_858_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_868_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_874_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_881_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_887_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_897_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_903_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_910_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_916_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_926_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_932_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_939_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_945_wire : std_logic_vector(0 downto 0);
    signal MUX_1007_wire : std_logic_vector(2 downto 0);
    signal MUX_1008_wire : std_logic_vector(2 downto 0);
    signal MUX_1009_wire : std_logic_vector(2 downto 0);
    signal MUX_1010_wire : std_logic_vector(2 downto 0);
    signal MUX_1034_wire : std_logic_vector(1 downto 0);
    signal MUX_1035_wire : std_logic_vector(1 downto 0);
    signal MUX_1036_wire : std_logic_vector(1 downto 0);
    signal MUX_1037_wire : std_logic_vector(1 downto 0);
    signal MUX_842_wire : std_logic_vector(0 downto 0);
    signal MUX_848_wire : std_logic_vector(0 downto 0);
    signal MUX_855_wire : std_logic_vector(0 downto 0);
    signal MUX_861_wire : std_logic_vector(0 downto 0);
    signal MUX_871_wire : std_logic_vector(0 downto 0);
    signal MUX_877_wire : std_logic_vector(0 downto 0);
    signal MUX_884_wire : std_logic_vector(0 downto 0);
    signal MUX_890_wire : std_logic_vector(0 downto 0);
    signal MUX_900_wire : std_logic_vector(0 downto 0);
    signal MUX_906_wire : std_logic_vector(0 downto 0);
    signal MUX_913_wire : std_logic_vector(0 downto 0);
    signal MUX_919_wire : std_logic_vector(0 downto 0);
    signal MUX_929_wire : std_logic_vector(0 downto 0);
    signal MUX_935_wire : std_logic_vector(0 downto 0);
    signal MUX_942_wire : std_logic_vector(0 downto 0);
    signal MUX_948_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1015_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_974_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_849_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_862_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_878_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_891_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_907_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_920_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_936_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_949_wire : std_logic_vector(0 downto 0);
    signal R_ZERO_1_977_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_1_983_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_1_991_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_1_999_wire_constant : std_logic_vector(0 downto 0);
    signal d0_835 : std_logic_vector(0 downto 0);
    signal konst_1001_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1004_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1006_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1019_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1023_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1027_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1031_wire_constant : std_logic_vector(1 downto 0);
    signal konst_833_wire_constant : std_logic_vector(7 downto 0);
    signal konst_838_wire_constant : std_logic_vector(1 downto 0);
    signal konst_841_wire_constant : std_logic_vector(0 downto 0);
    signal konst_844_wire_constant : std_logic_vector(1 downto 0);
    signal konst_847_wire_constant : std_logic_vector(0 downto 0);
    signal konst_851_wire_constant : std_logic_vector(1 downto 0);
    signal konst_854_wire_constant : std_logic_vector(0 downto 0);
    signal konst_857_wire_constant : std_logic_vector(1 downto 0);
    signal konst_860_wire_constant : std_logic_vector(0 downto 0);
    signal konst_867_wire_constant : std_logic_vector(1 downto 0);
    signal konst_870_wire_constant : std_logic_vector(0 downto 0);
    signal konst_873_wire_constant : std_logic_vector(1 downto 0);
    signal konst_876_wire_constant : std_logic_vector(0 downto 0);
    signal konst_880_wire_constant : std_logic_vector(1 downto 0);
    signal konst_883_wire_constant : std_logic_vector(0 downto 0);
    signal konst_886_wire_constant : std_logic_vector(1 downto 0);
    signal konst_889_wire_constant : std_logic_vector(0 downto 0);
    signal konst_896_wire_constant : std_logic_vector(1 downto 0);
    signal konst_899_wire_constant : std_logic_vector(0 downto 0);
    signal konst_902_wire_constant : std_logic_vector(1 downto 0);
    signal konst_905_wire_constant : std_logic_vector(0 downto 0);
    signal konst_909_wire_constant : std_logic_vector(1 downto 0);
    signal konst_912_wire_constant : std_logic_vector(0 downto 0);
    signal konst_915_wire_constant : std_logic_vector(1 downto 0);
    signal konst_918_wire_constant : std_logic_vector(0 downto 0);
    signal konst_925_wire_constant : std_logic_vector(1 downto 0);
    signal konst_928_wire_constant : std_logic_vector(0 downto 0);
    signal konst_931_wire_constant : std_logic_vector(1 downto 0);
    signal konst_934_wire_constant : std_logic_vector(0 downto 0);
    signal konst_938_wire_constant : std_logic_vector(1 downto 0);
    signal konst_941_wire_constant : std_logic_vector(0 downto 0);
    signal konst_944_wire_constant : std_logic_vector(1 downto 0);
    signal konst_947_wire_constant : std_logic_vector(0 downto 0);
    signal konst_980_wire_constant : std_logic_vector(2 downto 0);
    signal konst_985_wire_constant : std_logic_vector(1 downto 0);
    signal konst_988_wire_constant : std_logic_vector(2 downto 0);
    signal konst_993_wire_constant : std_logic_vector(1 downto 0);
    signal konst_996_wire_constant : std_logic_vector(2 downto 0);
    signal priority_1_validity_864 : std_logic_vector(0 downto 0);
    signal priority_2_validity_893 : std_logic_vector(0 downto 0);
    signal priority_3_validity_922 : std_logic_vector(0 downto 0);
    signal priority_4_validity_951 : std_logic_vector(0 downto 0);
    signal select_first_priority_956 : std_logic_vector(0 downto 0);
    signal select_fourth_priority_971 : std_logic_vector(0 downto 0);
    signal select_second_priority_961 : std_logic_vector(0 downto 0);
    signal select_third_priority_966 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_ZERO_1_977_wire_constant <= "0";
    R_ZERO_1_983_wire_constant <= "0";
    R_ZERO_1_991_wire_constant <= "0";
    R_ZERO_1_999_wire_constant <= "0";
    konst_1001_wire_constant <= "11";
    konst_1004_wire_constant <= "001";
    konst_1006_wire_constant <= "000";
    konst_1019_wire_constant <= "01";
    konst_1023_wire_constant <= "10";
    konst_1027_wire_constant <= "11";
    konst_1031_wire_constant <= "00";
    konst_833_wire_constant <= "00000000";
    konst_838_wire_constant <= "00";
    konst_841_wire_constant <= "0";
    konst_844_wire_constant <= "01";
    konst_847_wire_constant <= "0";
    konst_851_wire_constant <= "10";
    konst_854_wire_constant <= "0";
    konst_857_wire_constant <= "11";
    konst_860_wire_constant <= "0";
    konst_867_wire_constant <= "00";
    konst_870_wire_constant <= "0";
    konst_873_wire_constant <= "01";
    konst_876_wire_constant <= "0";
    konst_880_wire_constant <= "10";
    konst_883_wire_constant <= "0";
    konst_886_wire_constant <= "11";
    konst_889_wire_constant <= "0";
    konst_896_wire_constant <= "00";
    konst_899_wire_constant <= "0";
    konst_902_wire_constant <= "01";
    konst_905_wire_constant <= "0";
    konst_909_wire_constant <= "10";
    konst_912_wire_constant <= "0";
    konst_915_wire_constant <= "11";
    konst_918_wire_constant <= "0";
    konst_925_wire_constant <= "00";
    konst_928_wire_constant <= "0";
    konst_931_wire_constant <= "01";
    konst_934_wire_constant <= "0";
    konst_938_wire_constant <= "10";
    konst_941_wire_constant <= "0";
    konst_944_wire_constant <= "11";
    konst_947_wire_constant <= "0";
    konst_980_wire_constant <= "001";
    konst_985_wire_constant <= "01";
    konst_988_wire_constant <= "001";
    konst_993_wire_constant <= "10";
    konst_996_wire_constant <= "001";
    -- flow-through select operator MUX_1007_inst
    MUX_1007_wire <= ADD_u3_u3_1005_wire when (select_fourth_priority_971(0) /=  '0') else konst_1006_wire_constant;
    -- flow-through select operator MUX_1008_inst
    MUX_1008_wire <= ADD_u3_u3_997_wire when (select_third_priority_966(0) /=  '0') else MUX_1007_wire;
    -- flow-through select operator MUX_1009_inst
    MUX_1009_wire <= ADD_u3_u3_989_wire when (select_second_priority_961(0) /=  '0') else MUX_1008_wire;
    -- flow-through select operator MUX_1010_inst
    MUX_1010_wire <= ADD_u3_u3_981_wire when (select_first_priority_956(0) /=  '0') else MUX_1009_wire;
    -- flow-through select operator MUX_1011_inst
    next_active_packet_buffer <= active_packet_buffer when (NOT_u1_u1_974_wire(0) /=  '0') else MUX_1010_wire;
    -- flow-through select operator MUX_1034_inst
    MUX_1034_wire <= ADD_u2_u2_1032_wire when (select_fourth_priority_971(0) /=  '0') else priority_index_buffer;
    -- flow-through select operator MUX_1035_inst
    MUX_1035_wire <= ADD_u2_u2_1028_wire when (select_third_priority_966(0) /=  '0') else MUX_1034_wire;
    -- flow-through select operator MUX_1036_inst
    MUX_1036_wire <= ADD_u2_u2_1024_wire when (select_second_priority_961(0) /=  '0') else MUX_1035_wire;
    -- flow-through select operator MUX_1037_inst
    MUX_1037_wire <= ADD_u2_u2_1020_wire when (select_first_priority_956(0) /=  '0') else MUX_1036_wire;
    -- flow-through select operator MUX_1038_inst
    next_priority_index_buffer <= priority_index_buffer when (NOT_u1_u1_1015_wire(0) /=  '0') else MUX_1037_wire;
    -- flow-through select operator MUX_842_inst
    MUX_842_wire <= p1_valid_buffer when (EQ_u2_u1_839_wire(0) /=  '0') else konst_841_wire_constant;
    -- flow-through select operator MUX_848_inst
    MUX_848_wire <= p2_valid_buffer when (EQ_u2_u1_845_wire(0) /=  '0') else konst_847_wire_constant;
    -- flow-through select operator MUX_855_inst
    MUX_855_wire <= p3_valid_buffer when (EQ_u2_u1_852_wire(0) /=  '0') else konst_854_wire_constant;
    -- flow-through select operator MUX_861_inst
    MUX_861_wire <= p4_valid_buffer when (EQ_u2_u1_858_wire(0) /=  '0') else konst_860_wire_constant;
    -- flow-through select operator MUX_871_inst
    MUX_871_wire <= p2_valid_buffer when (EQ_u2_u1_868_wire(0) /=  '0') else konst_870_wire_constant;
    -- flow-through select operator MUX_877_inst
    MUX_877_wire <= p3_valid_buffer when (EQ_u2_u1_874_wire(0) /=  '0') else konst_876_wire_constant;
    -- flow-through select operator MUX_884_inst
    MUX_884_wire <= p4_valid_buffer when (EQ_u2_u1_881_wire(0) /=  '0') else konst_883_wire_constant;
    -- flow-through select operator MUX_890_inst
    MUX_890_wire <= p1_valid_buffer when (EQ_u2_u1_887_wire(0) /=  '0') else konst_889_wire_constant;
    -- flow-through select operator MUX_900_inst
    MUX_900_wire <= p3_valid_buffer when (EQ_u2_u1_897_wire(0) /=  '0') else konst_899_wire_constant;
    -- flow-through select operator MUX_906_inst
    MUX_906_wire <= p4_valid_buffer when (EQ_u2_u1_903_wire(0) /=  '0') else konst_905_wire_constant;
    -- flow-through select operator MUX_913_inst
    MUX_913_wire <= p1_valid_buffer when (EQ_u2_u1_910_wire(0) /=  '0') else konst_912_wire_constant;
    -- flow-through select operator MUX_919_inst
    MUX_919_wire <= p2_valid_buffer when (EQ_u2_u1_916_wire(0) /=  '0') else konst_918_wire_constant;
    -- flow-through select operator MUX_929_inst
    MUX_929_wire <= p4_valid_buffer when (EQ_u2_u1_926_wire(0) /=  '0') else konst_928_wire_constant;
    -- flow-through select operator MUX_935_inst
    MUX_935_wire <= p1_valid_buffer when (EQ_u2_u1_932_wire(0) /=  '0') else konst_934_wire_constant;
    -- flow-through select operator MUX_942_inst
    MUX_942_wire <= p2_valid_buffer when (EQ_u2_u1_939_wire(0) /=  '0') else konst_941_wire_constant;
    -- flow-through select operator MUX_948_inst
    MUX_948_wire <= p3_valid_buffer when (EQ_u2_u1_945_wire(0) /=  '0') else konst_947_wire_constant;
    -- flow through binary operator ADD_u2_u2_1002_inst
    ADD_u2_u2_1002_wire <= std_logic_vector(unsigned(priority_index_buffer) + unsigned(konst_1001_wire_constant));
    -- flow through binary operator ADD_u2_u2_1020_inst
    ADD_u2_u2_1020_wire <= std_logic_vector(unsigned(priority_index_buffer) + unsigned(konst_1019_wire_constant));
    -- flow through binary operator ADD_u2_u2_1024_inst
    ADD_u2_u2_1024_wire <= std_logic_vector(unsigned(priority_index_buffer) + unsigned(konst_1023_wire_constant));
    -- flow through binary operator ADD_u2_u2_1028_inst
    ADD_u2_u2_1028_wire <= std_logic_vector(unsigned(priority_index_buffer) + unsigned(konst_1027_wire_constant));
    -- flow through binary operator ADD_u2_u2_1032_inst
    ADD_u2_u2_1032_wire <= std_logic_vector(unsigned(priority_index_buffer) + unsigned(konst_1031_wire_constant));
    -- flow through binary operator ADD_u2_u2_986_inst
    ADD_u2_u2_986_wire <= std_logic_vector(unsigned(priority_index_buffer) + unsigned(konst_985_wire_constant));
    -- flow through binary operator ADD_u2_u2_994_inst
    ADD_u2_u2_994_wire <= std_logic_vector(unsigned(priority_index_buffer) + unsigned(konst_993_wire_constant));
    -- flow through binary operator ADD_u3_u3_1005_inst
    ADD_u3_u3_1005_wire <= std_logic_vector(unsigned(CONCAT_u1_u3_1003_wire) + unsigned(konst_1004_wire_constant));
    -- flow through binary operator ADD_u3_u3_981_inst
    ADD_u3_u3_981_wire <= std_logic_vector(unsigned(CONCAT_u1_u3_979_wire) + unsigned(konst_980_wire_constant));
    -- flow through binary operator ADD_u3_u3_989_inst
    ADD_u3_u3_989_wire <= std_logic_vector(unsigned(CONCAT_u1_u3_987_wire) + unsigned(konst_988_wire_constant));
    -- flow through binary operator ADD_u3_u3_997_inst
    ADD_u3_u3_997_wire <= std_logic_vector(unsigned(CONCAT_u1_u3_995_wire) + unsigned(konst_996_wire_constant));
    -- flow through binary operator AND_u1_u1_955_inst
    select_first_priority_956 <= (d0_835 and priority_1_validity_864);
    -- flow through binary operator AND_u1_u1_960_inst
    select_second_priority_961 <= (d0_835 and priority_2_validity_893);
    -- flow through binary operator AND_u1_u1_965_inst
    select_third_priority_966 <= (d0_835 and priority_3_validity_922);
    -- flow through binary operator AND_u1_u1_970_inst
    select_fourth_priority_971 <= (d0_835 and priority_4_validity_951);
    -- flow through binary operator CONCAT_u1_u3_1003_inst
    process(R_ZERO_1_999_wire_constant, ADD_u2_u2_1002_wire) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ZERO_1_999_wire_constant, ADD_u2_u2_1002_wire, tmp_var);
      CONCAT_u1_u3_1003_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u3_979_inst
    process(R_ZERO_1_977_wire_constant, priority_index_buffer) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ZERO_1_977_wire_constant, priority_index_buffer, tmp_var);
      CONCAT_u1_u3_979_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u3_987_inst
    process(R_ZERO_1_983_wire_constant, ADD_u2_u2_986_wire) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ZERO_1_983_wire_constant, ADD_u2_u2_986_wire, tmp_var);
      CONCAT_u1_u3_987_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u3_995_inst
    process(R_ZERO_1_991_wire_constant, ADD_u2_u2_994_wire) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ZERO_1_991_wire_constant, ADD_u2_u2_994_wire, tmp_var);
      CONCAT_u1_u3_995_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u2_u1_839_inst
    process(priority_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(priority_index_buffer, konst_838_wire_constant, tmp_var);
      EQ_u2_u1_839_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u2_u1_845_inst
    process(priority_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(priority_index_buffer, konst_844_wire_constant, tmp_var);
      EQ_u2_u1_845_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u2_u1_852_inst
    process(priority_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(priority_index_buffer, konst_851_wire_constant, tmp_var);
      EQ_u2_u1_852_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u2_u1_858_inst
    process(priority_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(priority_index_buffer, konst_857_wire_constant, tmp_var);
      EQ_u2_u1_858_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u2_u1_868_inst
    process(priority_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(priority_index_buffer, konst_867_wire_constant, tmp_var);
      EQ_u2_u1_868_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u2_u1_874_inst
    process(priority_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(priority_index_buffer, konst_873_wire_constant, tmp_var);
      EQ_u2_u1_874_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u2_u1_881_inst
    process(priority_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(priority_index_buffer, konst_880_wire_constant, tmp_var);
      EQ_u2_u1_881_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u2_u1_887_inst
    process(priority_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(priority_index_buffer, konst_886_wire_constant, tmp_var);
      EQ_u2_u1_887_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u2_u1_897_inst
    process(priority_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(priority_index_buffer, konst_896_wire_constant, tmp_var);
      EQ_u2_u1_897_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u2_u1_903_inst
    process(priority_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(priority_index_buffer, konst_902_wire_constant, tmp_var);
      EQ_u2_u1_903_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u2_u1_910_inst
    process(priority_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(priority_index_buffer, konst_909_wire_constant, tmp_var);
      EQ_u2_u1_910_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u2_u1_916_inst
    process(priority_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(priority_index_buffer, konst_915_wire_constant, tmp_var);
      EQ_u2_u1_916_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u2_u1_926_inst
    process(priority_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(priority_index_buffer, konst_925_wire_constant, tmp_var);
      EQ_u2_u1_926_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u2_u1_932_inst
    process(priority_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(priority_index_buffer, konst_931_wire_constant, tmp_var);
      EQ_u2_u1_932_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u2_u1_939_inst
    process(priority_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(priority_index_buffer, konst_938_wire_constant, tmp_var);
      EQ_u2_u1_939_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u2_u1_945_inst
    process(priority_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(priority_index_buffer, konst_944_wire_constant, tmp_var);
      EQ_u2_u1_945_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u8_u1_834_inst
    process(down_counter_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(down_counter_buffer, konst_833_wire_constant, tmp_var);
      d0_835 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1015_inst
    process(d0_835) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", d0_835, tmp_var);
      NOT_u1_u1_1015_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_974_inst
    process(d0_835) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", d0_835, tmp_var);
      NOT_u1_u1_974_wire <= tmp_var; -- 
    end process;
    -- flow through binary operator OR_u1_u1_849_inst
    OR_u1_u1_849_wire <= (MUX_842_wire or MUX_848_wire);
    -- flow through binary operator OR_u1_u1_862_inst
    OR_u1_u1_862_wire <= (MUX_855_wire or MUX_861_wire);
    -- flow through binary operator OR_u1_u1_863_inst
    priority_1_validity_864 <= (OR_u1_u1_849_wire or OR_u1_u1_862_wire);
    -- flow through binary operator OR_u1_u1_878_inst
    OR_u1_u1_878_wire <= (MUX_871_wire or MUX_877_wire);
    -- flow through binary operator OR_u1_u1_891_inst
    OR_u1_u1_891_wire <= (MUX_884_wire or MUX_890_wire);
    -- flow through binary operator OR_u1_u1_892_inst
    priority_2_validity_893 <= (OR_u1_u1_878_wire or OR_u1_u1_891_wire);
    -- flow through binary operator OR_u1_u1_907_inst
    OR_u1_u1_907_wire <= (MUX_900_wire or MUX_906_wire);
    -- flow through binary operator OR_u1_u1_920_inst
    OR_u1_u1_920_wire <= (MUX_913_wire or MUX_919_wire);
    -- flow through binary operator OR_u1_u1_921_inst
    priority_3_validity_922 <= (OR_u1_u1_907_wire or OR_u1_u1_920_wire);
    -- flow through binary operator OR_u1_u1_936_inst
    OR_u1_u1_936_wire <= (MUX_929_wire or MUX_935_wire);
    -- flow through binary operator OR_u1_u1_949_inst
    OR_u1_u1_949_wire <= (MUX_942_wire or MUX_948_wire);
    -- flow through binary operator OR_u1_u1_950_inst
    priority_4_validity_951 <= (OR_u1_u1_936_wire or OR_u1_u1_949_wire);
    -- 
  end Block; -- data_path
  -- 
end prioritySelect_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity updateCounter is -- 
  generic (tag_length : integer); 
  port ( -- 
    input_port : in  std_logic_vector(7 downto 0);
    output_port : in  std_logic_vector(7 downto 0);
    up : in  std_logic_vector(0 downto 0);
    continue : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(3 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(1 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(1 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity updateCounter;
architecture updateCounter_arch of updateCounter is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 17)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal input_port_buffer :  std_logic_vector(7 downto 0);
  signal input_port_update_enable: Boolean;
  signal output_port_buffer :  std_logic_vector(7 downto 0);
  signal output_port_update_enable: Boolean;
  signal up_buffer :  std_logic_vector(0 downto 0);
  signal up_update_enable: Boolean;
  -- output port buffer signals
  signal continue_buffer :  std_logic_vector(0 downto 0);
  signal continue_update_enable: Boolean;
  signal updateCounter_CP_294_start: Boolean;
  signal updateCounter_CP_294_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal array_obj_ref_177_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_177_index_sum_1_req_0 : boolean;
  signal array_obj_ref_177_store_0_ack_1 : boolean;
  signal array_obj_ref_177_store_0_req_1 : boolean;
  signal array_obj_ref_162_index_0_scale_req_1 : boolean;
  signal array_obj_ref_162_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_125_index_0_scale_req_0 : boolean;
  signal array_obj_ref_125_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_125_index_0_scale_req_1 : boolean;
  signal array_obj_ref_125_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_125_index_sum_1_req_0 : boolean;
  signal array_obj_ref_125_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_125_index_sum_1_req_1 : boolean;
  signal array_obj_ref_125_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_125_load_0_req_0 : boolean;
  signal array_obj_ref_125_load_0_ack_0 : boolean;
  signal array_obj_ref_177_store_0_ack_0 : boolean;
  signal array_obj_ref_125_load_0_req_1 : boolean;
  signal array_obj_ref_125_load_0_ack_1 : boolean;
  signal array_obj_ref_137_index_0_scale_req_0 : boolean;
  signal array_obj_ref_137_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_137_index_0_scale_req_1 : boolean;
  signal array_obj_ref_137_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_137_index_sum_1_req_0 : boolean;
  signal array_obj_ref_137_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_137_index_sum_1_req_1 : boolean;
  signal array_obj_ref_137_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_177_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_177_store_0_req_0 : boolean;
  signal array_obj_ref_137_load_0_req_0 : boolean;
  signal array_obj_ref_137_load_0_ack_0 : boolean;
  signal array_obj_ref_137_load_0_req_1 : boolean;
  signal array_obj_ref_137_load_0_ack_1 : boolean;
  signal array_obj_ref_177_index_0_scale_req_1 : boolean;
  signal array_obj_ref_150_index_0_scale_req_0 : boolean;
  signal array_obj_ref_150_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_177_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_150_index_0_scale_req_1 : boolean;
  signal array_obj_ref_150_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_150_index_sum_1_req_0 : boolean;
  signal array_obj_ref_150_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_177_index_sum_1_req_1 : boolean;
  signal array_obj_ref_150_index_sum_1_req_1 : boolean;
  signal array_obj_ref_150_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_150_load_0_req_0 : boolean;
  signal array_obj_ref_150_load_0_ack_0 : boolean;
  signal array_obj_ref_150_load_0_req_1 : boolean;
  signal array_obj_ref_150_load_0_ack_1 : boolean;
  signal array_obj_ref_162_index_0_scale_req_0 : boolean;
  signal array_obj_ref_162_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_162_index_sum_1_req_0 : boolean;
  signal array_obj_ref_162_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_162_index_sum_1_req_1 : boolean;
  signal array_obj_ref_162_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_162_load_0_req_0 : boolean;
  signal array_obj_ref_162_load_0_ack_0 : boolean;
  signal array_obj_ref_162_load_0_req_1 : boolean;
  signal array_obj_ref_162_load_0_ack_1 : boolean;
  signal array_obj_ref_185_index_0_scale_req_0 : boolean;
  signal array_obj_ref_185_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_185_index_0_scale_req_1 : boolean;
  signal array_obj_ref_185_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_185_index_sum_1_req_0 : boolean;
  signal array_obj_ref_185_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_185_index_sum_1_req_1 : boolean;
  signal array_obj_ref_185_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_185_load_0_req_0 : boolean;
  signal array_obj_ref_185_load_0_ack_0 : boolean;
  signal array_obj_ref_185_load_0_req_1 : boolean;
  signal array_obj_ref_185_load_0_ack_1 : boolean;
  signal array_obj_ref_197_index_0_scale_req_0 : boolean;
  signal array_obj_ref_197_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_197_index_0_scale_req_1 : boolean;
  signal array_obj_ref_197_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_197_index_sum_1_req_0 : boolean;
  signal array_obj_ref_197_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_197_index_sum_1_req_1 : boolean;
  signal array_obj_ref_197_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_197_load_0_req_0 : boolean;
  signal array_obj_ref_197_load_0_ack_0 : boolean;
  signal array_obj_ref_197_load_0_req_1 : boolean;
  signal array_obj_ref_197_load_0_ack_1 : boolean;
  signal array_obj_ref_207_index_0_scale_req_0 : boolean;
  signal array_obj_ref_207_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_207_index_0_scale_req_1 : boolean;
  signal array_obj_ref_207_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_207_index_sum_1_req_0 : boolean;
  signal array_obj_ref_207_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_207_index_sum_1_req_1 : boolean;
  signal array_obj_ref_207_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_207_load_0_req_0 : boolean;
  signal array_obj_ref_207_load_0_ack_0 : boolean;
  signal array_obj_ref_207_load_0_req_1 : boolean;
  signal array_obj_ref_207_load_0_ack_1 : boolean;
  signal OR_u2_u2_210_inst_req_0 : boolean;
  signal OR_u2_u2_210_inst_ack_0 : boolean;
  signal OR_u2_u2_210_inst_req_1 : boolean;
  signal OR_u2_u2_210_inst_ack_1 : boolean;
  signal array_obj_ref_177_index_0_scale_req_0 : boolean;
  signal array_obj_ref_177_index_0_scale_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "updateCounter_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 17) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= input_port;
  input_port_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(15 downto 8) <= output_port;
  output_port_buffer <= in_buffer_data_out(15 downto 8);
  in_buffer_data_in(16 downto 16) <= up;
  up_buffer <= in_buffer_data_out(16 downto 16);
  in_buffer_data_in(tag_length + 16 downto 17) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 16 downto 17);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  updateCounter_CP_294_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "updateCounter_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(0 downto 0) <= continue_buffer;
  continue <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= updateCounter_CP_294_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= updateCounter_CP_294_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= updateCounter_CP_294_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  updateCounter_CP_294: Block -- control-path 
    signal updateCounter_CP_294_elements: BooleanArray(68 downto 0);
    -- 
  begin -- 
    updateCounter_CP_294_elements(0) <= updateCounter_CP_294_start;
    updateCounter_CP_294_symbol <= updateCounter_CP_294_elements(68);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	15 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	14 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	10 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	34 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	43 
    -- CP-element group 0: 	36 
    -- CP-element group 0: 	46 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	37 
    -- CP-element group 0: 	38 
    -- CP-element group 0: 	39 
    -- CP-element group 0: 	41 
    -- CP-element group 0: 	60 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	58 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	54 
    -- CP-element group 0: 	55 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	45 
    -- CP-element group 0: 	50 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	17 
    -- CP-element group 0: 	19 
    -- CP-element group 0: 	30 
    -- CP-element group 0: 	31 
    -- CP-element group 0: 	21 
    -- CP-element group 0: 	22 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	26 
    -- CP-element group 0:  members (253) 
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_partial_sum_1_Update/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_partial_sum_1_update_start
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_scale_0_Update/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_scale_0_Update/cr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_resized_1
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_computed_1
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_partial_sum_1_update_start
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_update_start_
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_resized_0
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_computed_0
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_resize_0/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_resize_0/$exit
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_resize_0/index_resize_req
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_resize_0/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_scale_0_sample_start
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_scale_0_update_start
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_scale_0_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_scale_0_Sample/rr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_scale_0_Update/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_scale_0_Update/cr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_resized_1
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_computed_1
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_partial_sum_1_update_start
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_partial_sum_1_Update/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_partial_sum_1_Update/cr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_Update/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_Update/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_update_start_
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_resized_0
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_computed_0
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_resize_0/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_resize_0/$exit
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_resize_0/index_resize_req
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_resize_0/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_computed_1
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_scale_0_sample_start
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_scale_0_update_start
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_scale_0_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_scale_0_Sample/rr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_scale_0_Update/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_scale_0_Update/cr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_resized_1
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_computed_1
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_resized_1
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_partial_sum_1_update_start
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_partial_sum_1_Update/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_partial_sum_1_Update/cr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_Update/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_update_start_
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_resized_0
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_computed_0
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_resize_0/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_resize_0/$exit
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_resize_0/index_resize_req
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_resize_0/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_scale_0_Update/cr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_scale_0_sample_start
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_scale_0_update_start
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_scale_0_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_scale_0_Sample/rr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_scale_0_Update/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_scale_0_Update/cr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_resized_1
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_computed_1
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_scale_0_Update/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_partial_sum_1_update_start
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_partial_sum_1_Update/cr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_partial_sum_1_Update/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_partial_sum_1_Update/cr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_Update/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_update_start_
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_resized_0
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_computed_0
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_resize_0/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_resize_0/$exit
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_resize_0/index_resize_req
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_resize_0/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_scale_0_sample_start
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_scale_0_update_start
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_scale_0_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_scale_0_Sample/rr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_partial_sum_1_Update/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_partial_sum_1_Update/cr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_Update/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/OR_u2_u2_210_update_start_
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_update_start_
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_resized_0
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_computed_0
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_resize_0/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_resize_0/$exit
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_resize_0/index_resize_req
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_resize_0/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_scale_0_sample_start
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_scale_0_update_start
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_scale_0_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_scale_0_Sample/rr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_scale_0_Update/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_scale_0_Update/cr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_resized_1
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_computed_1
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_partial_sum_1_update_start
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_partial_sum_1_Update/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_partial_sum_1_Update/cr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_Update/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_update_start_
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_resized_0
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_computed_0
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_resize_0/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_resize_0/$exit
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_resize_0/index_resize_req
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_resize_0/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_scale_0_sample_start
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_scale_0_update_start
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_scale_0_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_scale_0_Sample/rr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_scale_0_Update/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_scale_0_Update/cr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_resized_1
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_computed_1
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_partial_sum_1_update_start
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_partial_sum_1_Update/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_partial_sum_1_Update/cr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_Update/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_update_start_
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_resized_0
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_computed_0
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_resize_0/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_resize_0/$exit
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_resize_0/index_resize_req
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_resize_0/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_scale_0_sample_start
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_scale_0_update_start
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_scale_0_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_scale_0_Sample/rr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_scale_0_Update/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_scale_0_Update/cr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_resized_1
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_computed_1
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_partial_sum_1_update_start
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_partial_sum_1_Update/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_partial_sum_1_Update/cr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_Update/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/OR_u2_u2_210_Update/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/OR_u2_u2_210_Update/cr
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_update_start_
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_resized_0
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_computed_0
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_resize_0/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_resize_0/$exit
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_resize_0/index_resize_req
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_resize_0/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_scale_0_sample_start
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_scale_0_update_start
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_scale_0_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_scale_0_Sample/rr
      -- 
    cr_391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_125_load_0_req_1); -- 
    rr_322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_125_index_0_scale_req_0); -- 
    cr_327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_125_index_0_scale_req_1); -- 
    cr_489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_137_load_0_req_1); -- 
    rr_420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_137_index_0_scale_req_0); -- 
    cr_587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_150_load_0_req_1); -- 
    rr_518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_150_index_0_scale_req_0); -- 
    cr_523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_150_index_0_scale_req_1); -- 
    cr_425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_137_index_0_scale_req_1); -- 
    cr_452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_137_index_sum_1_req_1); -- 
    cr_354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_125_index_sum_1_req_1); -- 
    cr_750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_185_index_sum_1_req_1); -- 
    cr_983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_207_load_0_req_1); -- 
    cr_946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_207_index_sum_1_req_1); -- 
    cr_885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_197_load_0_req_1); -- 
    rr_816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_197_index_0_scale_req_0); -- 
    cr_821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_197_index_0_scale_req_1); -- 
    cr_848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_197_index_sum_1_req_1); -- 
    cr_1054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_177_index_sum_1_req_1); -- 
    cr_1096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_177_store_0_req_1); -- 
    rr_1022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_177_index_0_scale_req_0); -- 
    cr_1027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_177_index_0_scale_req_1); -- 
    rr_914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_207_index_0_scale_req_0); -- 
    cr_919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_207_index_0_scale_req_1); -- 
    cr_550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_150_index_sum_1_req_1); -- 
    cr_998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => OR_u2_u2_210_inst_req_1); -- 
    cr_787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_185_load_0_req_1); -- 
    rr_718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_185_index_0_scale_req_0); -- 
    cr_723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_185_index_0_scale_req_1); -- 
    cr_685_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_685_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_162_load_0_req_1); -- 
    rr_616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_162_index_0_scale_req_0); -- 
    cr_621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_162_index_0_scale_req_1); -- 
    cr_648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(0), ack => array_obj_ref_162_index_sum_1_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	68 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_scale_0_sample_complete
      -- CP-element group 1: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_scale_0_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_scale_0_Sample/ra
      -- 
    ra_323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_125_index_0_scale_ack_0, ack => updateCounter_CP_294_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (4) 
      -- CP-element group 2: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_scaled_0
      -- CP-element group 2: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_scale_0_update_complete
      -- CP-element group 2: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_scale_0_Update/$exit
      -- CP-element group 2: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_index_scale_0_Update/ca
      -- 
    ca_328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_125_index_0_scale_ack_1, ack => updateCounter_CP_294_elements(2)); -- 
    -- CP-element group 3:  join  transition  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_partial_sum_1_sample_start
      -- CP-element group 3: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_partial_sum_1_Sample/$entry
      -- CP-element group 3: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_partial_sum_1_Sample/rr
      -- 
    rr_349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(3), ack => array_obj_ref_125_index_sum_1_req_0); -- 
    updateCounter_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "updateCounter_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= updateCounter_CP_294_elements(0) & updateCounter_CP_294_elements(2);
      gj_updateCounter_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => updateCounter_CP_294_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	68 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_partial_sum_1_sample_complete
      -- CP-element group 4: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_partial_sum_1_Sample/$exit
      -- CP-element group 4: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_partial_sum_1_Sample/ra
      -- 
    ra_350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_125_index_sum_1_ack_0, ack => updateCounter_CP_294_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (23) 
      -- CP-element group 5: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_sample_start_
      -- CP-element group 5: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_word_address_calculated
      -- CP-element group 5: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_root_address_calculated
      -- CP-element group 5: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_offset_calculated
      -- CP-element group 5: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_partial_sum_1_update_complete
      -- CP-element group 5: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_partial_sum_1_Update/$exit
      -- CP-element group 5: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_partial_sum_1_Update/ca
      -- CP-element group 5: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_final_index_sum_regn/$entry
      -- CP-element group 5: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_final_index_sum_regn/$exit
      -- CP-element group 5: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_final_index_sum_regn/req
      -- CP-element group 5: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_final_index_sum_regn/ack
      -- CP-element group 5: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_base_plus_offset/$entry
      -- CP-element group 5: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_base_plus_offset/$exit
      -- CP-element group 5: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_base_plus_offset/sum_rename_req
      -- CP-element group 5: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_base_plus_offset/sum_rename_ack
      -- CP-element group 5: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_word_addrgen/$entry
      -- CP-element group 5: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_word_addrgen/$exit
      -- CP-element group 5: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_word_addrgen/root_register_req
      -- CP-element group 5: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_word_addrgen/root_register_ack
      -- CP-element group 5: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_Sample/$entry
      -- CP-element group 5: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_Sample/word_access_start/$entry
      -- CP-element group 5: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_Sample/word_access_start/word_0/$entry
      -- CP-element group 5: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_Sample/word_access_start/word_0/rr
      -- 
    ca_355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_125_index_sum_1_ack_1, ack => updateCounter_CP_294_elements(5)); -- 
    rr_380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(5), ack => array_obj_ref_125_load_0_req_0); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	61 
    -- CP-element group 6:  members (5) 
      -- CP-element group 6: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_sample_completed_
      -- CP-element group 6: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_Sample/$exit
      -- CP-element group 6: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_Sample/word_access_start/$exit
      -- CP-element group 6: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_Sample/word_access_start/word_0/$exit
      -- CP-element group 6: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_Sample/word_access_start/word_0/ra
      -- 
    ra_381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_125_load_0_ack_0, ack => updateCounter_CP_294_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	29 
    -- CP-element group 7:  members (9) 
      -- CP-element group 7: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_update_completed_
      -- CP-element group 7: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_Update/$exit
      -- CP-element group 7: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_Update/word_access_complete/$exit
      -- CP-element group 7: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_Update/word_access_complete/word_0/$exit
      -- CP-element group 7: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_Update/word_access_complete/word_0/ca
      -- CP-element group 7: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_Update/array_obj_ref_125_Merge/$entry
      -- CP-element group 7: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_Update/array_obj_ref_125_Merge/$exit
      -- CP-element group 7: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_Update/array_obj_ref_125_Merge/merge_req
      -- CP-element group 7: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_Update/array_obj_ref_125_Merge/merge_ack
      -- 
    ca_392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_125_load_0_ack_1, ack => updateCounter_CP_294_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	68 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_scale_0_sample_complete
      -- CP-element group 8: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_scale_0_Sample/$exit
      -- CP-element group 8: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_scale_0_Sample/ra
      -- 
    ra_421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_137_index_0_scale_ack_0, ack => updateCounter_CP_294_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_scaled_0
      -- CP-element group 9: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_scale_0_update_complete
      -- CP-element group 9: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_scale_0_Update/$exit
      -- CP-element group 9: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_index_scale_0_Update/ca
      -- 
    ca_426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_137_index_0_scale_ack_1, ack => updateCounter_CP_294_elements(9)); -- 
    -- CP-element group 10:  join  transition  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	0 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_partial_sum_1_sample_start
      -- CP-element group 10: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_partial_sum_1_Sample/$entry
      -- CP-element group 10: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_partial_sum_1_Sample/rr
      -- 
    rr_447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(10), ack => array_obj_ref_137_index_sum_1_req_0); -- 
    updateCounter_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "updateCounter_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= updateCounter_CP_294_elements(0) & updateCounter_CP_294_elements(9);
      gj_updateCounter_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => updateCounter_CP_294_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	68 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_partial_sum_1_sample_complete
      -- CP-element group 11: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_partial_sum_1_Sample/$exit
      -- CP-element group 11: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_partial_sum_1_Sample/ra
      -- 
    ra_448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_137_index_sum_1_ack_0, ack => updateCounter_CP_294_elements(11)); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (23) 
      -- CP-element group 12: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_sample_start_
      -- CP-element group 12: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_word_address_calculated
      -- CP-element group 12: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_root_address_calculated
      -- CP-element group 12: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_offset_calculated
      -- CP-element group 12: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_partial_sum_1_update_complete
      -- CP-element group 12: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_partial_sum_1_Update/$exit
      -- CP-element group 12: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_partial_sum_1_Update/ca
      -- CP-element group 12: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_final_index_sum_regn/$entry
      -- CP-element group 12: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_final_index_sum_regn/$exit
      -- CP-element group 12: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_final_index_sum_regn/req
      -- CP-element group 12: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_final_index_sum_regn/ack
      -- CP-element group 12: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_base_plus_offset/$entry
      -- CP-element group 12: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_base_plus_offset/$exit
      -- CP-element group 12: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_base_plus_offset/sum_rename_req
      -- CP-element group 12: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_base_plus_offset/sum_rename_ack
      -- CP-element group 12: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_word_addrgen/$entry
      -- CP-element group 12: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_word_addrgen/$exit
      -- CP-element group 12: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_word_addrgen/root_register_req
      -- CP-element group 12: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_word_addrgen/root_register_ack
      -- CP-element group 12: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_Sample/$entry
      -- CP-element group 12: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_Sample/word_access_start/$entry
      -- CP-element group 12: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_Sample/word_access_start/word_0/$entry
      -- CP-element group 12: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_Sample/word_access_start/word_0/rr
      -- 
    ca_453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_137_index_sum_1_ack_1, ack => updateCounter_CP_294_elements(12)); -- 
    rr_478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(12), ack => array_obj_ref_137_load_0_req_0); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	62 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_sample_completed_
      -- CP-element group 13: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_Sample/$exit
      -- CP-element group 13: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_Sample/word_access_start/$exit
      -- CP-element group 13: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_Sample/word_access_start/word_0/ra
      -- 
    ra_479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_137_load_0_ack_0, ack => updateCounter_CP_294_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	0 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	29 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_update_completed_
      -- CP-element group 14: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_Update/$exit
      -- CP-element group 14: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_Update/word_access_complete/$exit
      -- CP-element group 14: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_Update/array_obj_ref_137_Merge/$entry
      -- CP-element group 14: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_Update/array_obj_ref_137_Merge/$exit
      -- CP-element group 14: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_Update/array_obj_ref_137_Merge/merge_req
      -- CP-element group 14: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_Update/array_obj_ref_137_Merge/merge_ack
      -- 
    ca_490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_137_load_0_ack_1, ack => updateCounter_CP_294_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	0 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	68 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_scale_0_sample_complete
      -- CP-element group 15: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_scale_0_Sample/$exit
      -- CP-element group 15: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_scale_0_Sample/ra
      -- 
    ra_519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_150_index_0_scale_ack_0, ack => updateCounter_CP_294_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (4) 
      -- CP-element group 16: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_scaled_0
      -- CP-element group 16: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_scale_0_update_complete
      -- CP-element group 16: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_scale_0_Update/$exit
      -- CP-element group 16: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_index_scale_0_Update/ca
      -- 
    ca_524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_150_index_0_scale_ack_1, ack => updateCounter_CP_294_elements(16)); -- 
    -- CP-element group 17:  join  transition  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	0 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_partial_sum_1_sample_start
      -- CP-element group 17: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_partial_sum_1_Sample/$entry
      -- CP-element group 17: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_partial_sum_1_Sample/rr
      -- 
    rr_545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(17), ack => array_obj_ref_150_index_sum_1_req_0); -- 
    updateCounter_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "updateCounter_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= updateCounter_CP_294_elements(0) & updateCounter_CP_294_elements(16);
      gj_updateCounter_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => updateCounter_CP_294_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	68 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_partial_sum_1_sample_complete
      -- CP-element group 18: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_partial_sum_1_Sample/$exit
      -- CP-element group 18: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_partial_sum_1_Sample/ra
      -- 
    ra_546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_150_index_sum_1_ack_0, ack => updateCounter_CP_294_elements(18)); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	0 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (23) 
      -- CP-element group 19: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_sample_start_
      -- CP-element group 19: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_word_address_calculated
      -- CP-element group 19: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_root_address_calculated
      -- CP-element group 19: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_offset_calculated
      -- CP-element group 19: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_partial_sum_1_update_complete
      -- CP-element group 19: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_partial_sum_1_Update/$exit
      -- CP-element group 19: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_partial_sum_1_Update/ca
      -- CP-element group 19: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_final_index_sum_regn/$entry
      -- CP-element group 19: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_final_index_sum_regn/$exit
      -- CP-element group 19: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_final_index_sum_regn/req
      -- CP-element group 19: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_final_index_sum_regn/ack
      -- CP-element group 19: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_base_plus_offset/$entry
      -- CP-element group 19: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_base_plus_offset/$exit
      -- CP-element group 19: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_base_plus_offset/sum_rename_req
      -- CP-element group 19: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_base_plus_offset/sum_rename_ack
      -- CP-element group 19: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_word_addrgen/$entry
      -- CP-element group 19: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_word_addrgen/$exit
      -- CP-element group 19: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_word_addrgen/root_register_req
      -- CP-element group 19: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_word_addrgen/root_register_ack
      -- CP-element group 19: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_Sample/$entry
      -- CP-element group 19: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_Sample/word_access_start/$entry
      -- CP-element group 19: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_Sample/word_access_start/word_0/$entry
      -- CP-element group 19: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_Sample/word_access_start/word_0/rr
      -- 
    ca_551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_150_index_sum_1_ack_1, ack => updateCounter_CP_294_elements(19)); -- 
    rr_576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(19), ack => array_obj_ref_150_load_0_req_0); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	63 
    -- CP-element group 20:  members (5) 
      -- CP-element group 20: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_sample_completed_
      -- CP-element group 20: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_Sample/$exit
      -- CP-element group 20: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_Sample/word_access_start/$exit
      -- CP-element group 20: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_Sample/word_access_start/word_0/$exit
      -- CP-element group 20: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_Sample/word_access_start/word_0/ra
      -- 
    ra_577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_150_load_0_ack_0, ack => updateCounter_CP_294_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	0 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	29 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_update_completed_
      -- CP-element group 21: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_Update/$exit
      -- CP-element group 21: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_Update/word_access_complete/$exit
      -- CP-element group 21: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_Update/word_access_complete/word_0/$exit
      -- CP-element group 21: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_Update/word_access_complete/word_0/ca
      -- CP-element group 21: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_Update/array_obj_ref_150_Merge/$entry
      -- CP-element group 21: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_Update/array_obj_ref_150_Merge/$exit
      -- CP-element group 21: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_Update/array_obj_ref_150_Merge/merge_req
      -- CP-element group 21: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_Update/array_obj_ref_150_Merge/merge_ack
      -- 
    ca_588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_150_load_0_ack_1, ack => updateCounter_CP_294_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	0 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	68 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_scale_0_sample_complete
      -- CP-element group 22: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_scale_0_Sample/$exit
      -- CP-element group 22: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_scale_0_Sample/ra
      -- 
    ra_617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_162_index_0_scale_ack_0, ack => updateCounter_CP_294_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (4) 
      -- CP-element group 23: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_scale_0_Update/$exit
      -- CP-element group 23: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_scale_0_Update/ca
      -- CP-element group 23: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_scaled_0
      -- CP-element group 23: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_index_scale_0_update_complete
      -- 
    ca_622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_162_index_0_scale_ack_1, ack => updateCounter_CP_294_elements(23)); -- 
    -- CP-element group 24:  join  transition  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_partial_sum_1_sample_start
      -- CP-element group 24: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_partial_sum_1_Sample/$entry
      -- CP-element group 24: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_partial_sum_1_Sample/rr
      -- 
    rr_643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(24), ack => array_obj_ref_162_index_sum_1_req_0); -- 
    updateCounter_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "updateCounter_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= updateCounter_CP_294_elements(0) & updateCounter_CP_294_elements(23);
      gj_updateCounter_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => updateCounter_CP_294_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	68 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_partial_sum_1_sample_complete
      -- CP-element group 25: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_partial_sum_1_Sample/$exit
      -- CP-element group 25: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_partial_sum_1_Sample/ra
      -- 
    ra_644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_162_index_sum_1_ack_0, ack => updateCounter_CP_294_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	0 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (23) 
      -- CP-element group 26: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_partial_sum_1_update_complete
      -- CP-element group 26: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_sample_start_
      -- CP-element group 26: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_word_address_calculated
      -- CP-element group 26: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_root_address_calculated
      -- CP-element group 26: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_offset_calculated
      -- CP-element group 26: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_partial_sum_1_Update/$exit
      -- CP-element group 26: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_partial_sum_1_Update/ca
      -- CP-element group 26: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_final_index_sum_regn/$entry
      -- CP-element group 26: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_final_index_sum_regn/$exit
      -- CP-element group 26: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_final_index_sum_regn/req
      -- CP-element group 26: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_final_index_sum_regn/ack
      -- CP-element group 26: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_base_plus_offset/$entry
      -- CP-element group 26: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_base_plus_offset/$exit
      -- CP-element group 26: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_base_plus_offset/sum_rename_req
      -- CP-element group 26: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_base_plus_offset/sum_rename_ack
      -- CP-element group 26: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_word_addrgen/$entry
      -- CP-element group 26: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_word_addrgen/$exit
      -- CP-element group 26: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_word_addrgen/root_register_req
      -- CP-element group 26: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_word_addrgen/root_register_ack
      -- CP-element group 26: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_Sample/$entry
      -- CP-element group 26: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_Sample/word_access_start/$entry
      -- CP-element group 26: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_Sample/word_access_start/word_0/$entry
      -- CP-element group 26: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_Sample/word_access_start/word_0/rr
      -- 
    ca_649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_162_index_sum_1_ack_1, ack => updateCounter_CP_294_elements(26)); -- 
    rr_674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(26), ack => array_obj_ref_162_load_0_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	64 
    -- CP-element group 27:  members (5) 
      -- CP-element group 27: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_sample_completed_
      -- CP-element group 27: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_Sample/$exit
      -- CP-element group 27: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_Sample/word_access_start/$exit
      -- CP-element group 27: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_Sample/word_access_start/word_0/$exit
      -- CP-element group 27: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_Sample/word_access_start/word_0/ra
      -- 
    ra_675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_162_load_0_ack_0, ack => updateCounter_CP_294_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (9) 
      -- CP-element group 28: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_update_completed_
      -- CP-element group 28: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_Update/$exit
      -- CP-element group 28: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_Update/word_access_complete/$exit
      -- CP-element group 28: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_Update/word_access_complete/word_0/$exit
      -- CP-element group 28: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_Update/word_access_complete/word_0/ca
      -- CP-element group 28: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_Update/array_obj_ref_162_Merge/$entry
      -- CP-element group 28: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_Update/array_obj_ref_162_Merge/$exit
      -- CP-element group 28: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_Update/array_obj_ref_162_Merge/merge_req
      -- CP-element group 28: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_Update/array_obj_ref_162_Merge/merge_ack
      -- 
    ca_686_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_162_load_0_ack_1, ack => updateCounter_CP_294_elements(28)); -- 
    -- CP-element group 29:  join  transition  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	7 
    -- CP-element group 29: 	14 
    -- CP-element group 29: 	28 
    -- CP-element group 29: 	43 
    -- CP-element group 29: 	36 
    -- CP-element group 29: 	50 
    -- CP-element group 29: 	21 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	51 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 assign_stmt_121_to_assign_stmt_211/OR_u2_u2_210_sample_start_
      -- CP-element group 29: 	 assign_stmt_121_to_assign_stmt_211/OR_u2_u2_210_Sample/$entry
      -- CP-element group 29: 	 assign_stmt_121_to_assign_stmt_211/OR_u2_u2_210_Sample/rr
      -- 
    rr_993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(29), ack => OR_u2_u2_210_inst_req_0); -- 
    updateCounter_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 33) := "updateCounter_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= updateCounter_CP_294_elements(7) & updateCounter_CP_294_elements(14) & updateCounter_CP_294_elements(28) & updateCounter_CP_294_elements(43) & updateCounter_CP_294_elements(36) & updateCounter_CP_294_elements(50) & updateCounter_CP_294_elements(21);
      gj_updateCounter_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => updateCounter_CP_294_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	0 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	68 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_scale_0_sample_complete
      -- CP-element group 30: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_scale_0_Sample/$exit
      -- CP-element group 30: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_scale_0_Sample/ra
      -- 
    ra_719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_185_index_0_scale_ack_0, ack => updateCounter_CP_294_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	0 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_scaled_0
      -- CP-element group 31: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_scale_0_update_complete
      -- CP-element group 31: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_scale_0_Update/$exit
      -- CP-element group 31: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_index_scale_0_Update/ca
      -- 
    ca_724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_185_index_0_scale_ack_1, ack => updateCounter_CP_294_elements(31)); -- 
    -- CP-element group 32:  join  transition  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_partial_sum_1_sample_start
      -- CP-element group 32: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_partial_sum_1_Sample/$entry
      -- CP-element group 32: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_partial_sum_1_Sample/rr
      -- 
    rr_745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(32), ack => array_obj_ref_185_index_sum_1_req_0); -- 
    updateCounter_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "updateCounter_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= updateCounter_CP_294_elements(0) & updateCounter_CP_294_elements(31);
      gj_updateCounter_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => updateCounter_CP_294_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	68 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_partial_sum_1_sample_complete
      -- CP-element group 33: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_partial_sum_1_Sample/$exit
      -- CP-element group 33: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_partial_sum_1_Sample/ra
      -- 
    ra_746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_185_index_sum_1_ack_0, ack => updateCounter_CP_294_elements(33)); -- 
    -- CP-element group 34:  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	0 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (23) 
      -- CP-element group 34: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_sample_start_
      -- CP-element group 34: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_word_address_calculated
      -- CP-element group 34: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_root_address_calculated
      -- CP-element group 34: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_offset_calculated
      -- CP-element group 34: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_partial_sum_1_update_complete
      -- CP-element group 34: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_partial_sum_1_Update/$exit
      -- CP-element group 34: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_partial_sum_1_Update/ca
      -- CP-element group 34: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_final_index_sum_regn/$entry
      -- CP-element group 34: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_final_index_sum_regn/$exit
      -- CP-element group 34: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_final_index_sum_regn/req
      -- CP-element group 34: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_final_index_sum_regn/ack
      -- CP-element group 34: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_base_plus_offset/$entry
      -- CP-element group 34: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_base_plus_offset/$exit
      -- CP-element group 34: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_base_plus_offset/sum_rename_req
      -- CP-element group 34: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_base_plus_offset/sum_rename_ack
      -- CP-element group 34: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_word_addrgen/$entry
      -- CP-element group 34: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_word_addrgen/$exit
      -- CP-element group 34: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_word_addrgen/root_register_req
      -- CP-element group 34: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_word_addrgen/root_register_ack
      -- CP-element group 34: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_Sample/$entry
      -- CP-element group 34: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_Sample/word_access_start/$entry
      -- CP-element group 34: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_Sample/word_access_start/word_0/$entry
      -- CP-element group 34: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_Sample/word_access_start/word_0/rr
      -- 
    ca_751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_185_index_sum_1_ack_1, ack => updateCounter_CP_294_elements(34)); -- 
    rr_776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(34), ack => array_obj_ref_185_load_0_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	65 
    -- CP-element group 35:  members (5) 
      -- CP-element group 35: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_sample_completed_
      -- CP-element group 35: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_Sample/$exit
      -- CP-element group 35: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_Sample/word_access_start/$exit
      -- CP-element group 35: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_Sample/word_access_start/word_0/$exit
      -- CP-element group 35: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_Sample/word_access_start/word_0/ra
      -- 
    ra_777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_185_load_0_ack_0, ack => updateCounter_CP_294_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	29 
    -- CP-element group 36:  members (9) 
      -- CP-element group 36: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_update_completed_
      -- CP-element group 36: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_Update/$exit
      -- CP-element group 36: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_Update/word_access_complete/$exit
      -- CP-element group 36: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_Update/word_access_complete/word_0/$exit
      -- CP-element group 36: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_Update/word_access_complete/word_0/ca
      -- CP-element group 36: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_Update/array_obj_ref_185_Merge/$entry
      -- CP-element group 36: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_Update/array_obj_ref_185_Merge/$exit
      -- CP-element group 36: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_Update/array_obj_ref_185_Merge/merge_req
      -- CP-element group 36: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_Update/array_obj_ref_185_Merge/merge_ack
      -- 
    ca_788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_185_load_0_ack_1, ack => updateCounter_CP_294_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	0 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	68 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_scale_0_sample_complete
      -- CP-element group 37: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_scale_0_Sample/$exit
      -- CP-element group 37: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_scale_0_Sample/ra
      -- 
    ra_817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_197_index_0_scale_ack_0, ack => updateCounter_CP_294_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	0 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_scaled_0
      -- CP-element group 38: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_scale_0_update_complete
      -- CP-element group 38: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_scale_0_Update/$exit
      -- CP-element group 38: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_index_scale_0_Update/ca
      -- 
    ca_822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_197_index_0_scale_ack_1, ack => updateCounter_CP_294_elements(38)); -- 
    -- CP-element group 39:  join  transition  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	0 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_partial_sum_1_sample_start
      -- CP-element group 39: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_partial_sum_1_Sample/$entry
      -- CP-element group 39: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_partial_sum_1_Sample/rr
      -- 
    rr_843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(39), ack => array_obj_ref_197_index_sum_1_req_0); -- 
    updateCounter_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "updateCounter_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= updateCounter_CP_294_elements(0) & updateCounter_CP_294_elements(38);
      gj_updateCounter_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => updateCounter_CP_294_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	68 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_partial_sum_1_sample_complete
      -- CP-element group 40: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_partial_sum_1_Sample/$exit
      -- CP-element group 40: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_partial_sum_1_Sample/ra
      -- 
    ra_844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_197_index_sum_1_ack_0, ack => updateCounter_CP_294_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	0 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (23) 
      -- CP-element group 41: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_sample_start_
      -- CP-element group 41: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_word_address_calculated
      -- CP-element group 41: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_root_address_calculated
      -- CP-element group 41: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_offset_calculated
      -- CP-element group 41: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_partial_sum_1_update_complete
      -- CP-element group 41: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_partial_sum_1_Update/$exit
      -- CP-element group 41: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_partial_sum_1_Update/ca
      -- CP-element group 41: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_final_index_sum_regn/$entry
      -- CP-element group 41: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_final_index_sum_regn/$exit
      -- CP-element group 41: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_final_index_sum_regn/req
      -- CP-element group 41: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_final_index_sum_regn/ack
      -- CP-element group 41: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_base_plus_offset/$entry
      -- CP-element group 41: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_base_plus_offset/$exit
      -- CP-element group 41: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_base_plus_offset/sum_rename_req
      -- CP-element group 41: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_base_plus_offset/sum_rename_ack
      -- CP-element group 41: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_word_addrgen/$entry
      -- CP-element group 41: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_word_addrgen/$exit
      -- CP-element group 41: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_word_addrgen/root_register_req
      -- CP-element group 41: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_word_addrgen/root_register_ack
      -- CP-element group 41: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_Sample/$entry
      -- CP-element group 41: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_Sample/word_access_start/$entry
      -- CP-element group 41: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_Sample/word_access_start/word_0/$entry
      -- CP-element group 41: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_Sample/word_access_start/word_0/rr
      -- 
    ca_849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_197_index_sum_1_ack_1, ack => updateCounter_CP_294_elements(41)); -- 
    rr_874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(41), ack => array_obj_ref_197_load_0_req_0); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	66 
    -- CP-element group 42:  members (5) 
      -- CP-element group 42: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_sample_completed_
      -- CP-element group 42: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_Sample/$exit
      -- CP-element group 42: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_Sample/word_access_start/$exit
      -- CP-element group 42: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_Sample/word_access_start/word_0/$exit
      -- CP-element group 42: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_Sample/word_access_start/word_0/ra
      -- 
    ra_875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_197_load_0_ack_0, ack => updateCounter_CP_294_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	0 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	29 
    -- CP-element group 43:  members (9) 
      -- CP-element group 43: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_update_completed_
      -- CP-element group 43: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_Update/$exit
      -- CP-element group 43: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_Update/word_access_complete/$exit
      -- CP-element group 43: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_Update/word_access_complete/word_0/$exit
      -- CP-element group 43: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_Update/word_access_complete/word_0/ca
      -- CP-element group 43: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_Update/array_obj_ref_197_Merge/$entry
      -- CP-element group 43: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_Update/array_obj_ref_197_Merge/$exit
      -- CP-element group 43: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_Update/array_obj_ref_197_Merge/merge_req
      -- CP-element group 43: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_Update/array_obj_ref_197_Merge/merge_ack
      -- 
    ca_886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_197_load_0_ack_1, ack => updateCounter_CP_294_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	68 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_scale_0_sample_complete
      -- CP-element group 44: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_scale_0_Sample/$exit
      -- CP-element group 44: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_scale_0_Sample/ra
      -- 
    ra_915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_207_index_0_scale_ack_0, ack => updateCounter_CP_294_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	0 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_scaled_0
      -- CP-element group 45: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_scale_0_update_complete
      -- CP-element group 45: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_scale_0_Update/$exit
      -- CP-element group 45: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_index_scale_0_Update/ca
      -- 
    ca_920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_207_index_0_scale_ack_1, ack => updateCounter_CP_294_elements(45)); -- 
    -- CP-element group 46:  join  transition  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	0 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_partial_sum_1_sample_start
      -- CP-element group 46: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_partial_sum_1_Sample/$entry
      -- CP-element group 46: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_partial_sum_1_Sample/rr
      -- 
    rr_941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(46), ack => array_obj_ref_207_index_sum_1_req_0); -- 
    updateCounter_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "updateCounter_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= updateCounter_CP_294_elements(0) & updateCounter_CP_294_elements(45);
      gj_updateCounter_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => updateCounter_CP_294_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	68 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_partial_sum_1_sample_complete
      -- CP-element group 47: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_partial_sum_1_Sample/$exit
      -- CP-element group 47: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_partial_sum_1_Sample/ra
      -- 
    ra_942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_207_index_sum_1_ack_0, ack => updateCounter_CP_294_elements(47)); -- 
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (23) 
      -- CP-element group 48: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_sample_start_
      -- CP-element group 48: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_word_address_calculated
      -- CP-element group 48: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_root_address_calculated
      -- CP-element group 48: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_offset_calculated
      -- CP-element group 48: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_partial_sum_1_update_complete
      -- CP-element group 48: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_partial_sum_1_Update/$exit
      -- CP-element group 48: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_partial_sum_1_Update/ca
      -- CP-element group 48: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_final_index_sum_regn/$entry
      -- CP-element group 48: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_final_index_sum_regn/$exit
      -- CP-element group 48: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_final_index_sum_regn/req
      -- CP-element group 48: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_final_index_sum_regn/ack
      -- CP-element group 48: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_base_plus_offset/$entry
      -- CP-element group 48: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_base_plus_offset/$exit
      -- CP-element group 48: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_base_plus_offset/sum_rename_req
      -- CP-element group 48: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_base_plus_offset/sum_rename_ack
      -- CP-element group 48: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_word_addrgen/$entry
      -- CP-element group 48: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_word_addrgen/$exit
      -- CP-element group 48: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_word_addrgen/root_register_req
      -- CP-element group 48: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_word_addrgen/root_register_ack
      -- CP-element group 48: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_Sample/$entry
      -- CP-element group 48: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_Sample/word_access_start/$entry
      -- CP-element group 48: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_Sample/word_access_start/word_0/$entry
      -- CP-element group 48: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_Sample/word_access_start/word_0/rr
      -- 
    ca_947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_207_index_sum_1_ack_1, ack => updateCounter_CP_294_elements(48)); -- 
    rr_972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(48), ack => array_obj_ref_207_load_0_req_0); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	67 
    -- CP-element group 49:  members (5) 
      -- CP-element group 49: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_sample_completed_
      -- CP-element group 49: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_Sample/$exit
      -- CP-element group 49: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_Sample/word_access_start/$exit
      -- CP-element group 49: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_Sample/word_access_start/word_0/$exit
      -- CP-element group 49: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_Sample/word_access_start/word_0/ra
      -- 
    ra_973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_207_load_0_ack_0, ack => updateCounter_CP_294_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	0 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	29 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_update_completed_
      -- CP-element group 50: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_Update/$exit
      -- CP-element group 50: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_Update/word_access_complete/$exit
      -- CP-element group 50: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_Update/word_access_complete/word_0/$exit
      -- CP-element group 50: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_Update/word_access_complete/word_0/ca
      -- CP-element group 50: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_Update/array_obj_ref_207_Merge/$entry
      -- CP-element group 50: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_Update/array_obj_ref_207_Merge/$exit
      -- CP-element group 50: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_Update/array_obj_ref_207_Merge/merge_req
      -- CP-element group 50: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_Update/array_obj_ref_207_Merge/merge_ack
      -- 
    ca_984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_207_load_0_ack_1, ack => updateCounter_CP_294_elements(50)); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	29 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 assign_stmt_121_to_assign_stmt_211/OR_u2_u2_210_sample_completed_
      -- CP-element group 51: 	 assign_stmt_121_to_assign_stmt_211/OR_u2_u2_210_Sample/$exit
      -- CP-element group 51: 	 assign_stmt_121_to_assign_stmt_211/OR_u2_u2_210_Sample/ra
      -- 
    ra_994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u2_u2_210_inst_ack_0, ack => updateCounter_CP_294_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 assign_stmt_121_to_assign_stmt_211/OR_u2_u2_210_update_completed_
      -- CP-element group 52: 	 assign_stmt_121_to_assign_stmt_211/OR_u2_u2_210_Update/$exit
      -- CP-element group 52: 	 assign_stmt_121_to_assign_stmt_211/OR_u2_u2_210_Update/ca
      -- 
    ca_999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u2_u2_210_inst_ack_1, ack => updateCounter_CP_294_elements(52)); -- 
    -- CP-element group 53:  join  transition  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	61 
    -- CP-element group 53: 	58 
    -- CP-element group 53: 	52 
    -- CP-element group 53: 	62 
    -- CP-element group 53: 	63 
    -- CP-element group 53: 	64 
    -- CP-element group 53: 	65 
    -- CP-element group 53: 	66 
    -- CP-element group 53: 	67 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	59 
    -- CP-element group 53:  members (9) 
      -- CP-element group 53: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_Sample/word_access_start/word_0/$entry
      -- CP-element group 53: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_Sample/word_access_start/$entry
      -- CP-element group 53: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_Sample/array_obj_ref_177_Split/split_ack
      -- CP-element group 53: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_Sample/array_obj_ref_177_Split/split_req
      -- CP-element group 53: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_Sample/array_obj_ref_177_Split/$exit
      -- CP-element group 53: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_Sample/array_obj_ref_177_Split/$entry
      -- CP-element group 53: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_Sample/$entry
      -- CP-element group 53: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_Sample/word_access_start/word_0/rr
      -- CP-element group 53: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_sample_start_
      -- 
    rr_1085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(53), ack => array_obj_ref_177_store_0_req_0); -- 
    updateCounter_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 33) := "updateCounter_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= updateCounter_CP_294_elements(61) & updateCounter_CP_294_elements(58) & updateCounter_CP_294_elements(52) & updateCounter_CP_294_elements(62) & updateCounter_CP_294_elements(63) & updateCounter_CP_294_elements(64) & updateCounter_CP_294_elements(65) & updateCounter_CP_294_elements(66) & updateCounter_CP_294_elements(67);
      gj_updateCounter_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => updateCounter_CP_294_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	0 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	68 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_scale_0_sample_complete
      -- CP-element group 54: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_scale_0_Sample/$exit
      -- CP-element group 54: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_scale_0_Sample/ra
      -- 
    ra_1023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_177_index_0_scale_ack_0, ack => updateCounter_CP_294_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	0 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_scale_0_Update/ca
      -- CP-element group 55: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_scale_0_Update/$exit
      -- CP-element group 55: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_scaled_0
      -- CP-element group 55: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_index_scale_0_update_complete
      -- 
    ca_1028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_177_index_0_scale_ack_1, ack => updateCounter_CP_294_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_partial_sum_1_Sample/rr
      -- CP-element group 56: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_partial_sum_1_Sample/$entry
      -- CP-element group 56: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_partial_sum_1_sample_start
      -- 
    rr_1049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateCounter_CP_294_elements(56), ack => array_obj_ref_177_index_sum_1_req_0); -- 
    updateCounter_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "updateCounter_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= updateCounter_CP_294_elements(0) & updateCounter_CP_294_elements(55);
      gj_updateCounter_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => updateCounter_CP_294_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	68 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_partial_sum_1_Sample/ra
      -- CP-element group 57: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_partial_sum_1_Sample/$exit
      -- CP-element group 57: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_partial_sum_1_sample_complete
      -- 
    ra_1050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_177_index_sum_1_ack_0, ack => updateCounter_CP_294_elements(57)); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	0 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	53 
    -- CP-element group 58:  members (18) 
      -- CP-element group 58: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_partial_sum_1_Update/$exit
      -- CP-element group 58: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_partial_sum_1_update_complete
      -- CP-element group 58: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_word_addrgen/root_register_ack
      -- CP-element group 58: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_word_addrgen/root_register_req
      -- CP-element group 58: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_word_addrgen/$exit
      -- CP-element group 58: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_word_addrgen/$entry
      -- CP-element group 58: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_base_plus_offset/sum_rename_ack
      -- CP-element group 58: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_base_plus_offset/sum_rename_req
      -- CP-element group 58: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_base_plus_offset/$exit
      -- CP-element group 58: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_base_plus_offset/$entry
      -- CP-element group 58: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_final_index_sum_regn/ack
      -- CP-element group 58: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_final_index_sum_regn/req
      -- CP-element group 58: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_final_index_sum_regn/$exit
      -- CP-element group 58: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_final_index_sum_regn/$entry
      -- CP-element group 58: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_partial_sum_1_Update/ca
      -- CP-element group 58: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_word_address_calculated
      -- CP-element group 58: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_root_address_calculated
      -- CP-element group 58: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_offset_calculated
      -- 
    ca_1055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_177_index_sum_1_ack_1, ack => updateCounter_CP_294_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	53 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (5) 
      -- CP-element group 59: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_Sample/word_access_start/$exit
      -- CP-element group 59: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_Sample/$exit
      -- CP-element group 59: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_Sample/word_access_start/word_0/ra
      -- CP-element group 59: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_Sample/word_access_start/word_0/$exit
      -- CP-element group 59: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_sample_completed_
      -- 
    ra_1086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_177_store_0_ack_0, ack => updateCounter_CP_294_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	0 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	68 
    -- CP-element group 60:  members (5) 
      -- CP-element group 60: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_Update/word_access_complete/word_0/ca
      -- CP-element group 60: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_Update/word_access_complete/word_0/$exit
      -- CP-element group 60: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_Update/word_access_complete/$exit
      -- CP-element group 60: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_Update/$exit
      -- CP-element group 60: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_177_update_completed_
      -- 
    ca_1097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_177_store_0_ack_1, ack => updateCounter_CP_294_elements(60)); -- 
    -- CP-element group 61:  transition  delay-element  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	6 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	53 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_125_array_obj_ref_177_delay
      -- 
    -- Element group updateCounter_CP_294_elements(61) is a control-delay.
    cp_element_61_delay: control_delay_element  generic map(name => " 61_delay", delay_value => 1)  port map(req => updateCounter_CP_294_elements(6), ack => updateCounter_CP_294_elements(61), clk => clk, reset =>reset);
    -- CP-element group 62:  transition  delay-element  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	13 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	53 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_137_array_obj_ref_177_delay
      -- 
    -- Element group updateCounter_CP_294_elements(62) is a control-delay.
    cp_element_62_delay: control_delay_element  generic map(name => " 62_delay", delay_value => 1)  port map(req => updateCounter_CP_294_elements(13), ack => updateCounter_CP_294_elements(62), clk => clk, reset =>reset);
    -- CP-element group 63:  transition  delay-element  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	20 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	53 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_150_array_obj_ref_177_delay
      -- 
    -- Element group updateCounter_CP_294_elements(63) is a control-delay.
    cp_element_63_delay: control_delay_element  generic map(name => " 63_delay", delay_value => 1)  port map(req => updateCounter_CP_294_elements(20), ack => updateCounter_CP_294_elements(63), clk => clk, reset =>reset);
    -- CP-element group 64:  transition  delay-element  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	27 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	53 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_162_array_obj_ref_177_delay
      -- 
    -- Element group updateCounter_CP_294_elements(64) is a control-delay.
    cp_element_64_delay: control_delay_element  generic map(name => " 64_delay", delay_value => 1)  port map(req => updateCounter_CP_294_elements(27), ack => updateCounter_CP_294_elements(64), clk => clk, reset =>reset);
    -- CP-element group 65:  transition  delay-element  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	35 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	53 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_185_array_obj_ref_177_delay
      -- 
    -- Element group updateCounter_CP_294_elements(65) is a control-delay.
    cp_element_65_delay: control_delay_element  generic map(name => " 65_delay", delay_value => 1)  port map(req => updateCounter_CP_294_elements(35), ack => updateCounter_CP_294_elements(65), clk => clk, reset =>reset);
    -- CP-element group 66:  transition  delay-element  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	42 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	53 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_197_array_obj_ref_177_delay
      -- 
    -- Element group updateCounter_CP_294_elements(66) is a control-delay.
    cp_element_66_delay: control_delay_element  generic map(name => " 66_delay", delay_value => 1)  port map(req => updateCounter_CP_294_elements(42), ack => updateCounter_CP_294_elements(66), clk => clk, reset =>reset);
    -- CP-element group 67:  transition  delay-element  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	49 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	53 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 assign_stmt_121_to_assign_stmt_211/array_obj_ref_207_array_obj_ref_177_delay
      -- 
    -- Element group updateCounter_CP_294_elements(67) is a control-delay.
    cp_element_67_delay: control_delay_element  generic map(name => " 67_delay", delay_value => 1)  port map(req => updateCounter_CP_294_elements(49), ack => updateCounter_CP_294_elements(67), clk => clk, reset =>reset);
    -- CP-element group 68:  join  transition  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	1 
    -- CP-element group 68: 	15 
    -- CP-element group 68: 	8 
    -- CP-element group 68: 	11 
    -- CP-element group 68: 	4 
    -- CP-element group 68: 	33 
    -- CP-element group 68: 	47 
    -- CP-element group 68: 	37 
    -- CP-element group 68: 	40 
    -- CP-element group 68: 	60 
    -- CP-element group 68: 	57 
    -- CP-element group 68: 	54 
    -- CP-element group 68: 	44 
    -- CP-element group 68: 	18 
    -- CP-element group 68: 	30 
    -- CP-element group 68: 	22 
    -- CP-element group 68: 	25 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 $exit
      -- CP-element group 68: 	 assign_stmt_121_to_assign_stmt_211/$exit
      -- 
    updateCounter_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 33) := "updateCounter_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= updateCounter_CP_294_elements(1) & updateCounter_CP_294_elements(15) & updateCounter_CP_294_elements(8) & updateCounter_CP_294_elements(11) & updateCounter_CP_294_elements(4) & updateCounter_CP_294_elements(33) & updateCounter_CP_294_elements(47) & updateCounter_CP_294_elements(37) & updateCounter_CP_294_elements(40) & updateCounter_CP_294_elements(60) & updateCounter_CP_294_elements(57) & updateCounter_CP_294_elements(54) & updateCounter_CP_294_elements(44) & updateCounter_CP_294_elements(18) & updateCounter_CP_294_elements(30) & updateCounter_CP_294_elements(22) & updateCounter_CP_294_elements(25);
      gj_updateCounter_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => updateCounter_CP_294_elements(68), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u2_u2_199_wire : std_logic_vector(1 downto 0);
    signal AND_u1_u1_131_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_143_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_156_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_168_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_182_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_194_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_130_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_142_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_155_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_167_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_181_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_193_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_152_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_164_wire : std_logic_vector(0 downto 0);
    signal MUX_134_wire : std_logic_vector(0 downto 0);
    signal MUX_146_wire : std_logic_vector(0 downto 0);
    signal MUX_159_wire : std_logic_vector(0 downto 0);
    signal MUX_171_wire : std_logic_vector(0 downto 0);
    signal MUX_189_wire : std_logic_vector(1 downto 0);
    signal MUX_201_wire : std_logic_vector(1 downto 0);
    signal MUX_209_wire : std_logic_vector(1 downto 0);
    signal NOT_u1_u1_204_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_147_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_172_wire : std_logic_vector(0 downto 0);
    signal OR_u2_u2_202_wire : std_logic_vector(1 downto 0);
    signal OR_u2_u2_210_wire : std_logic_vector(1 downto 0);
    signal R_input_port_123_resized : std_logic_vector(3 downto 0);
    signal R_input_port_123_scaled : std_logic_vector(3 downto 0);
    signal R_input_port_135_resized : std_logic_vector(3 downto 0);
    signal R_input_port_135_scaled : std_logic_vector(3 downto 0);
    signal R_input_port_148_resized : std_logic_vector(3 downto 0);
    signal R_input_port_148_scaled : std_logic_vector(3 downto 0);
    signal R_input_port_160_resized : std_logic_vector(3 downto 0);
    signal R_input_port_160_scaled : std_logic_vector(3 downto 0);
    signal R_input_port_175_resized : std_logic_vector(3 downto 0);
    signal R_input_port_175_scaled : std_logic_vector(3 downto 0);
    signal R_input_port_183_resized : std_logic_vector(3 downto 0);
    signal R_input_port_183_scaled : std_logic_vector(3 downto 0);
    signal R_input_port_195_resized : std_logic_vector(3 downto 0);
    signal R_input_port_195_scaled : std_logic_vector(3 downto 0);
    signal R_input_port_205_resized : std_logic_vector(3 downto 0);
    signal R_input_port_205_scaled : std_logic_vector(3 downto 0);
    signal R_output_port_124_resized : std_logic_vector(3 downto 0);
    signal R_output_port_124_scaled : std_logic_vector(3 downto 0);
    signal R_output_port_136_resized : std_logic_vector(3 downto 0);
    signal R_output_port_136_scaled : std_logic_vector(3 downto 0);
    signal R_output_port_149_resized : std_logic_vector(3 downto 0);
    signal R_output_port_149_scaled : std_logic_vector(3 downto 0);
    signal R_output_port_161_resized : std_logic_vector(3 downto 0);
    signal R_output_port_161_scaled : std_logic_vector(3 downto 0);
    signal R_output_port_176_resized : std_logic_vector(3 downto 0);
    signal R_output_port_176_scaled : std_logic_vector(3 downto 0);
    signal R_output_port_184_resized : std_logic_vector(3 downto 0);
    signal R_output_port_184_scaled : std_logic_vector(3 downto 0);
    signal R_output_port_196_resized : std_logic_vector(3 downto 0);
    signal R_output_port_196_scaled : std_logic_vector(3 downto 0);
    signal R_output_port_206_resized : std_logic_vector(3 downto 0);
    signal R_output_port_206_scaled : std_logic_vector(3 downto 0);
    signal SUB_u2_u2_187_wire : std_logic_vector(1 downto 0);
    signal UGT_u2_u1_127_wire : std_logic_vector(0 downto 0);
    signal ULT_u2_u1_139_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_125_data_0 : std_logic_vector(1 downto 0);
    signal array_obj_ref_125_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_125_index_partial_sum_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_125_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_125_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_125_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_125_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_125_wire : std_logic_vector(1 downto 0);
    signal array_obj_ref_125_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_125_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_137_data_0 : std_logic_vector(1 downto 0);
    signal array_obj_ref_137_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_137_index_partial_sum_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_137_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_137_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_137_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_137_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_137_wire : std_logic_vector(1 downto 0);
    signal array_obj_ref_137_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_137_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_150_data_0 : std_logic_vector(1 downto 0);
    signal array_obj_ref_150_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_150_index_partial_sum_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_150_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_150_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_150_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_150_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_150_wire : std_logic_vector(1 downto 0);
    signal array_obj_ref_150_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_150_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_162_data_0 : std_logic_vector(1 downto 0);
    signal array_obj_ref_162_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_162_index_partial_sum_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_162_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_162_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_162_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_162_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_162_wire : std_logic_vector(1 downto 0);
    signal array_obj_ref_162_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_162_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_177_data_0 : std_logic_vector(1 downto 0);
    signal array_obj_ref_177_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_177_index_partial_sum_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_177_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_177_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_177_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_177_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_177_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_177_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_185_data_0 : std_logic_vector(1 downto 0);
    signal array_obj_ref_185_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_185_index_partial_sum_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_185_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_185_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_185_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_185_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_185_wire : std_logic_vector(1 downto 0);
    signal array_obj_ref_185_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_185_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_197_data_0 : std_logic_vector(1 downto 0);
    signal array_obj_ref_197_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_197_index_partial_sum_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_197_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_197_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_197_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_197_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_197_wire : std_logic_vector(1 downto 0);
    signal array_obj_ref_197_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_197_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_207_data_0 : std_logic_vector(1 downto 0);
    signal array_obj_ref_207_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_207_index_partial_sum_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_207_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_207_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_207_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_207_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_207_wire : std_logic_vector(1 downto 0);
    signal array_obj_ref_207_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_207_word_offset_0 : std_logic_vector(3 downto 0);
    signal down_121 : std_logic_vector(0 downto 0);
    signal konst_126_wire_constant : std_logic_vector(1 downto 0);
    signal konst_129_wire_constant : std_logic_vector(0 downto 0);
    signal konst_132_wire_constant : std_logic_vector(0 downto 0);
    signal konst_133_wire_constant : std_logic_vector(0 downto 0);
    signal konst_138_wire_constant : std_logic_vector(1 downto 0);
    signal konst_141_wire_constant : std_logic_vector(0 downto 0);
    signal konst_144_wire_constant : std_logic_vector(0 downto 0);
    signal konst_145_wire_constant : std_logic_vector(0 downto 0);
    signal konst_151_wire_constant : std_logic_vector(1 downto 0);
    signal konst_154_wire_constant : std_logic_vector(0 downto 0);
    signal konst_157_wire_constant : std_logic_vector(0 downto 0);
    signal konst_158_wire_constant : std_logic_vector(0 downto 0);
    signal konst_163_wire_constant : std_logic_vector(1 downto 0);
    signal konst_166_wire_constant : std_logic_vector(0 downto 0);
    signal konst_169_wire_constant : std_logic_vector(0 downto 0);
    signal konst_170_wire_constant : std_logic_vector(0 downto 0);
    signal konst_180_wire_constant : std_logic_vector(0 downto 0);
    signal konst_186_wire_constant : std_logic_vector(1 downto 0);
    signal konst_188_wire_constant : std_logic_vector(1 downto 0);
    signal konst_192_wire_constant : std_logic_vector(0 downto 0);
    signal konst_198_wire_constant : std_logic_vector(1 downto 0);
    signal konst_200_wire_constant : std_logic_vector(1 downto 0);
    signal konst_208_wire_constant : std_logic_vector(1 downto 0);
    -- 
  begin -- 
    array_obj_ref_125_offset_scale_factor_0 <= "0100";
    array_obj_ref_125_offset_scale_factor_1 <= "0001";
    array_obj_ref_125_resized_base_address <= "0000";
    array_obj_ref_125_word_offset_0 <= "0000";
    array_obj_ref_137_offset_scale_factor_0 <= "0100";
    array_obj_ref_137_offset_scale_factor_1 <= "0001";
    array_obj_ref_137_resized_base_address <= "0000";
    array_obj_ref_137_word_offset_0 <= "0000";
    array_obj_ref_150_offset_scale_factor_0 <= "0100";
    array_obj_ref_150_offset_scale_factor_1 <= "0001";
    array_obj_ref_150_resized_base_address <= "0000";
    array_obj_ref_150_word_offset_0 <= "0000";
    array_obj_ref_162_offset_scale_factor_0 <= "0100";
    array_obj_ref_162_offset_scale_factor_1 <= "0001";
    array_obj_ref_162_resized_base_address <= "0000";
    array_obj_ref_162_word_offset_0 <= "0000";
    array_obj_ref_177_offset_scale_factor_0 <= "0100";
    array_obj_ref_177_offset_scale_factor_1 <= "0001";
    array_obj_ref_177_resized_base_address <= "0000";
    array_obj_ref_177_word_offset_0 <= "0000";
    array_obj_ref_185_offset_scale_factor_0 <= "0100";
    array_obj_ref_185_offset_scale_factor_1 <= "0001";
    array_obj_ref_185_resized_base_address <= "0000";
    array_obj_ref_185_word_offset_0 <= "0000";
    array_obj_ref_197_offset_scale_factor_0 <= "0100";
    array_obj_ref_197_offset_scale_factor_1 <= "0001";
    array_obj_ref_197_resized_base_address <= "0000";
    array_obj_ref_197_word_offset_0 <= "0000";
    array_obj_ref_207_offset_scale_factor_0 <= "0100";
    array_obj_ref_207_offset_scale_factor_1 <= "0001";
    array_obj_ref_207_resized_base_address <= "0000";
    array_obj_ref_207_word_offset_0 <= "0000";
    konst_126_wire_constant <= "11";
    konst_129_wire_constant <= "1";
    konst_132_wire_constant <= "1";
    konst_133_wire_constant <= "0";
    konst_138_wire_constant <= "01";
    konst_141_wire_constant <= "1";
    konst_144_wire_constant <= "1";
    konst_145_wire_constant <= "0";
    konst_151_wire_constant <= "00";
    konst_154_wire_constant <= "1";
    konst_157_wire_constant <= "0";
    konst_158_wire_constant <= "0";
    konst_163_wire_constant <= "00";
    konst_166_wire_constant <= "1";
    konst_169_wire_constant <= "0";
    konst_170_wire_constant <= "0";
    konst_180_wire_constant <= "1";
    konst_186_wire_constant <= "01";
    konst_188_wire_constant <= "00";
    konst_192_wire_constant <= "1";
    konst_198_wire_constant <= "01";
    konst_200_wire_constant <= "00";
    konst_208_wire_constant <= "00";
    -- flow-through select operator MUX_134_inst
    MUX_134_wire <= konst_132_wire_constant when (AND_u1_u1_131_wire(0) /=  '0') else konst_133_wire_constant;
    -- flow-through select operator MUX_146_inst
    MUX_146_wire <= konst_144_wire_constant when (AND_u1_u1_143_wire(0) /=  '0') else konst_145_wire_constant;
    -- flow-through select operator MUX_159_inst
    MUX_159_wire <= konst_157_wire_constant when (AND_u1_u1_156_wire(0) /=  '0') else konst_158_wire_constant;
    -- flow-through select operator MUX_171_inst
    MUX_171_wire <= konst_169_wire_constant when (AND_u1_u1_168_wire(0) /=  '0') else konst_170_wire_constant;
    -- flow-through select operator MUX_189_inst
    MUX_189_wire <= SUB_u2_u2_187_wire when (AND_u1_u1_182_wire(0) /=  '0') else konst_188_wire_constant;
    -- flow-through select operator MUX_201_inst
    MUX_201_wire <= ADD_u2_u2_199_wire when (AND_u1_u1_194_wire(0) /=  '0') else konst_200_wire_constant;
    -- flow-through select operator MUX_209_inst
    MUX_209_wire <= array_obj_ref_207_wire when (NOT_u1_u1_204_wire(0) /=  '0') else konst_208_wire_constant;
    -- equivalence array_obj_ref_125_addr_0
    process(array_obj_ref_125_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_125_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_125_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_125_gather_scatter
    process(array_obj_ref_125_data_0) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(1 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_125_data_0;
      ov(1 downto 0) := iv;
      array_obj_ref_125_wire <= ov(1 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_125_index_0_resize
    process(input_port_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := input_port_buffer;
      ov := iv(3 downto 0);
      R_input_port_123_resized <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_125_index_1_rename
    process(R_output_port_124_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_output_port_124_resized;
      ov(3 downto 0) := iv;
      R_output_port_124_scaled <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_125_index_1_resize
    process(output_port_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := output_port_buffer;
      ov := iv(3 downto 0);
      R_output_port_124_resized <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_125_index_offset
    process(array_obj_ref_125_index_partial_sum_1) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_125_index_partial_sum_1;
      ov(3 downto 0) := iv;
      array_obj_ref_125_final_offset <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_125_root_address_inst
    process(array_obj_ref_125_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_125_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_125_root_address <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_137_addr_0
    process(array_obj_ref_137_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_137_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_137_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_137_gather_scatter
    process(array_obj_ref_137_data_0) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(1 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_137_data_0;
      ov(1 downto 0) := iv;
      array_obj_ref_137_wire <= ov(1 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_137_index_0_resize
    process(input_port_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := input_port_buffer;
      ov := iv(3 downto 0);
      R_input_port_135_resized <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_137_index_1_rename
    process(R_output_port_136_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_output_port_136_resized;
      ov(3 downto 0) := iv;
      R_output_port_136_scaled <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_137_index_1_resize
    process(output_port_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := output_port_buffer;
      ov := iv(3 downto 0);
      R_output_port_136_resized <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_137_index_offset
    process(array_obj_ref_137_index_partial_sum_1) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_137_index_partial_sum_1;
      ov(3 downto 0) := iv;
      array_obj_ref_137_final_offset <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_137_root_address_inst
    process(array_obj_ref_137_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_137_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_137_root_address <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_150_addr_0
    process(array_obj_ref_150_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_150_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_150_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_150_gather_scatter
    process(array_obj_ref_150_data_0) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(1 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_150_data_0;
      ov(1 downto 0) := iv;
      array_obj_ref_150_wire <= ov(1 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_150_index_0_resize
    process(input_port_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := input_port_buffer;
      ov := iv(3 downto 0);
      R_input_port_148_resized <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_150_index_1_rename
    process(R_output_port_149_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_output_port_149_resized;
      ov(3 downto 0) := iv;
      R_output_port_149_scaled <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_150_index_1_resize
    process(output_port_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := output_port_buffer;
      ov := iv(3 downto 0);
      R_output_port_149_resized <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_150_index_offset
    process(array_obj_ref_150_index_partial_sum_1) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_150_index_partial_sum_1;
      ov(3 downto 0) := iv;
      array_obj_ref_150_final_offset <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_150_root_address_inst
    process(array_obj_ref_150_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_150_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_150_root_address <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_162_addr_0
    process(array_obj_ref_162_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_162_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_162_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_162_gather_scatter
    process(array_obj_ref_162_data_0) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(1 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_162_data_0;
      ov(1 downto 0) := iv;
      array_obj_ref_162_wire <= ov(1 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_162_index_0_resize
    process(input_port_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := input_port_buffer;
      ov := iv(3 downto 0);
      R_input_port_160_resized <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_162_index_1_rename
    process(R_output_port_161_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_output_port_161_resized;
      ov(3 downto 0) := iv;
      R_output_port_161_scaled <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_162_index_1_resize
    process(output_port_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := output_port_buffer;
      ov := iv(3 downto 0);
      R_output_port_161_resized <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_162_index_offset
    process(array_obj_ref_162_index_partial_sum_1) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_162_index_partial_sum_1;
      ov(3 downto 0) := iv;
      array_obj_ref_162_final_offset <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_162_root_address_inst
    process(array_obj_ref_162_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_162_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_162_root_address <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_177_addr_0
    process(array_obj_ref_177_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_177_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_177_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_177_gather_scatter
    process(OR_u2_u2_210_wire) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(1 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := OR_u2_u2_210_wire;
      ov(1 downto 0) := iv;
      array_obj_ref_177_data_0 <= ov(1 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_177_index_0_resize
    process(input_port_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := input_port_buffer;
      ov := iv(3 downto 0);
      R_input_port_175_resized <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_177_index_1_rename
    process(R_output_port_176_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_output_port_176_resized;
      ov(3 downto 0) := iv;
      R_output_port_176_scaled <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_177_index_1_resize
    process(output_port_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := output_port_buffer;
      ov := iv(3 downto 0);
      R_output_port_176_resized <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_177_index_offset
    process(array_obj_ref_177_index_partial_sum_1) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_177_index_partial_sum_1;
      ov(3 downto 0) := iv;
      array_obj_ref_177_final_offset <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_177_root_address_inst
    process(array_obj_ref_177_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_177_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_177_root_address <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_185_addr_0
    process(array_obj_ref_185_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_185_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_185_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_185_gather_scatter
    process(array_obj_ref_185_data_0) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(1 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_185_data_0;
      ov(1 downto 0) := iv;
      array_obj_ref_185_wire <= ov(1 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_185_index_0_resize
    process(input_port_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := input_port_buffer;
      ov := iv(3 downto 0);
      R_input_port_183_resized <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_185_index_1_rename
    process(R_output_port_184_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_output_port_184_resized;
      ov(3 downto 0) := iv;
      R_output_port_184_scaled <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_185_index_1_resize
    process(output_port_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := output_port_buffer;
      ov := iv(3 downto 0);
      R_output_port_184_resized <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_185_index_offset
    process(array_obj_ref_185_index_partial_sum_1) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_185_index_partial_sum_1;
      ov(3 downto 0) := iv;
      array_obj_ref_185_final_offset <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_185_root_address_inst
    process(array_obj_ref_185_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_185_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_185_root_address <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_197_addr_0
    process(array_obj_ref_197_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_197_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_197_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_197_gather_scatter
    process(array_obj_ref_197_data_0) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(1 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_197_data_0;
      ov(1 downto 0) := iv;
      array_obj_ref_197_wire <= ov(1 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_197_index_0_resize
    process(input_port_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := input_port_buffer;
      ov := iv(3 downto 0);
      R_input_port_195_resized <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_197_index_1_rename
    process(R_output_port_196_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_output_port_196_resized;
      ov(3 downto 0) := iv;
      R_output_port_196_scaled <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_197_index_1_resize
    process(output_port_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := output_port_buffer;
      ov := iv(3 downto 0);
      R_output_port_196_resized <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_197_index_offset
    process(array_obj_ref_197_index_partial_sum_1) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_197_index_partial_sum_1;
      ov(3 downto 0) := iv;
      array_obj_ref_197_final_offset <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_197_root_address_inst
    process(array_obj_ref_197_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_197_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_197_root_address <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_207_addr_0
    process(array_obj_ref_207_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_207_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_207_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_207_gather_scatter
    process(array_obj_ref_207_data_0) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(1 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_207_data_0;
      ov(1 downto 0) := iv;
      array_obj_ref_207_wire <= ov(1 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_207_index_0_resize
    process(input_port_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := input_port_buffer;
      ov := iv(3 downto 0);
      R_input_port_205_resized <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_207_index_1_rename
    process(R_output_port_206_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_output_port_206_resized;
      ov(3 downto 0) := iv;
      R_output_port_206_scaled <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_207_index_1_resize
    process(output_port_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := output_port_buffer;
      ov := iv(3 downto 0);
      R_output_port_206_resized <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_207_index_offset
    process(array_obj_ref_207_index_partial_sum_1) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_207_index_partial_sum_1;
      ov(3 downto 0) := iv;
      array_obj_ref_207_final_offset <= ov(3 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_207_root_address_inst
    process(array_obj_ref_207_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_207_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_207_root_address <= ov(3 downto 0);
      --
    end process;
    -- flow through binary operator ADD_u2_u2_199_inst
    ADD_u2_u2_199_wire <= std_logic_vector(unsigned(array_obj_ref_197_wire) + unsigned(konst_198_wire_constant));
    -- flow through binary operator AND_u1_u1_131_inst
    AND_u1_u1_131_wire <= (UGT_u2_u1_127_wire and EQ_u1_u1_130_wire);
    -- flow through binary operator AND_u1_u1_143_inst
    AND_u1_u1_143_wire <= (ULT_u2_u1_139_wire and EQ_u1_u1_142_wire);
    -- flow through binary operator AND_u1_u1_156_inst
    AND_u1_u1_156_wire <= (EQ_u2_u1_152_wire and EQ_u1_u1_155_wire);
    -- flow through binary operator AND_u1_u1_168_inst
    AND_u1_u1_168_wire <= (EQ_u2_u1_164_wire and EQ_u1_u1_167_wire);
    -- flow through binary operator AND_u1_u1_182_inst
    AND_u1_u1_182_wire <= (continue_buffer and EQ_u1_u1_181_wire);
    -- flow through binary operator AND_u1_u1_194_inst
    AND_u1_u1_194_wire <= (continue_buffer and EQ_u1_u1_193_wire);
    -- flow through binary operator EQ_u1_u1_130_inst
    process(down_121) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(down_121, konst_129_wire_constant, tmp_var);
      EQ_u1_u1_130_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u1_u1_142_inst
    process(up_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(up_buffer, konst_141_wire_constant, tmp_var);
      EQ_u1_u1_142_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u1_u1_155_inst
    process(up_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(up_buffer, konst_154_wire_constant, tmp_var);
      EQ_u1_u1_155_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u1_u1_167_inst
    process(down_121) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(down_121, konst_166_wire_constant, tmp_var);
      EQ_u1_u1_167_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u1_u1_181_inst
    process(down_121) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(down_121, konst_180_wire_constant, tmp_var);
      EQ_u1_u1_181_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u1_u1_193_inst
    process(up_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(up_buffer, konst_192_wire_constant, tmp_var);
      EQ_u1_u1_193_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u2_u1_152_inst
    process(array_obj_ref_150_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(array_obj_ref_150_wire, konst_151_wire_constant, tmp_var);
      EQ_u2_u1_152_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u2_u1_164_inst
    process(array_obj_ref_162_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(array_obj_ref_162_wire, konst_163_wire_constant, tmp_var);
      EQ_u2_u1_164_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_120_inst
    process(up_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", up_buffer, tmp_var);
      down_121 <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_204_inst
    process(continue_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", continue_buffer, tmp_var);
      NOT_u1_u1_204_wire <= tmp_var; -- 
    end process;
    -- flow through binary operator OR_u1_u1_147_inst
    OR_u1_u1_147_wire <= (MUX_134_wire or MUX_146_wire);
    -- flow through binary operator OR_u1_u1_172_inst
    OR_u1_u1_172_wire <= (MUX_159_wire or MUX_171_wire);
    -- flow through binary operator OR_u1_u1_173_inst
    continue_buffer <= (OR_u1_u1_147_wire or OR_u1_u1_172_wire);
    -- flow through binary operator OR_u2_u2_202_inst
    OR_u2_u2_202_wire <= (MUX_189_wire or MUX_201_wire);
    -- shared split operator group (21) : OR_u2_u2_210_inst 
    ApIntOr_group_21: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(1 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= OR_u2_u2_202_wire & MUX_209_wire;
      OR_u2_u2_210_wire <= data_out(1 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u2_u2_210_inst_req_0;
      OR_u2_u2_210_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u2_u2_210_inst_req_1;
      OR_u2_u2_210_inst_ack_1 <= ackR_unguarded(0);
      ApIntOr_group_21_gI: SplitGuardInterface generic map(name => "ApIntOr_group_21_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_21",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 2,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 2, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 2,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- flow through binary operator SUB_u2_u2_187_inst
    SUB_u2_u2_187_wire <= std_logic_vector(unsigned(array_obj_ref_185_wire) - unsigned(konst_186_wire_constant));
    -- flow through binary operator UGT_u2_u1_127_inst
    process(array_obj_ref_125_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(array_obj_ref_125_wire, konst_126_wire_constant, tmp_var);
      UGT_u2_u1_127_wire <= tmp_var; --
    end process;
    -- flow through binary operator ULT_u2_u1_139_inst
    process(array_obj_ref_137_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(array_obj_ref_137_wire, konst_138_wire_constant, tmp_var);
      ULT_u2_u1_139_wire <= tmp_var; --
    end process;
    -- shared split operator group (25) : array_obj_ref_125_index_0_scale array_obj_ref_137_index_0_scale array_obj_ref_150_index_0_scale array_obj_ref_162_index_0_scale array_obj_ref_185_index_0_scale array_obj_ref_197_index_0_scale array_obj_ref_207_index_0_scale array_obj_ref_177_index_0_scale 
    ApIntMul_group_25: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 7 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(7 downto 0) := (7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      data_in <= R_input_port_123_resized & R_input_port_135_resized & R_input_port_148_resized & R_input_port_160_resized & R_input_port_183_resized & R_input_port_195_resized & R_input_port_205_resized & R_input_port_175_resized;
      R_input_port_123_scaled <= data_out(31 downto 28);
      R_input_port_135_scaled <= data_out(27 downto 24);
      R_input_port_148_scaled <= data_out(23 downto 20);
      R_input_port_160_scaled <= data_out(19 downto 16);
      R_input_port_183_scaled <= data_out(15 downto 12);
      R_input_port_195_scaled <= data_out(11 downto 8);
      R_input_port_205_scaled <= data_out(7 downto 4);
      R_input_port_175_scaled <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      reqL_unguarded(7) <= array_obj_ref_125_index_0_scale_req_0;
      reqL_unguarded(6) <= array_obj_ref_137_index_0_scale_req_0;
      reqL_unguarded(5) <= array_obj_ref_150_index_0_scale_req_0;
      reqL_unguarded(4) <= array_obj_ref_162_index_0_scale_req_0;
      reqL_unguarded(3) <= array_obj_ref_185_index_0_scale_req_0;
      reqL_unguarded(2) <= array_obj_ref_197_index_0_scale_req_0;
      reqL_unguarded(1) <= array_obj_ref_207_index_0_scale_req_0;
      reqL_unguarded(0) <= array_obj_ref_177_index_0_scale_req_0;
      array_obj_ref_125_index_0_scale_ack_0 <= ackL_unguarded(7);
      array_obj_ref_137_index_0_scale_ack_0 <= ackL_unguarded(6);
      array_obj_ref_150_index_0_scale_ack_0 <= ackL_unguarded(5);
      array_obj_ref_162_index_0_scale_ack_0 <= ackL_unguarded(4);
      array_obj_ref_185_index_0_scale_ack_0 <= ackL_unguarded(3);
      array_obj_ref_197_index_0_scale_ack_0 <= ackL_unguarded(2);
      array_obj_ref_207_index_0_scale_ack_0 <= ackL_unguarded(1);
      array_obj_ref_177_index_0_scale_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(7) <= array_obj_ref_125_index_0_scale_req_1;
      reqR_unguarded(6) <= array_obj_ref_137_index_0_scale_req_1;
      reqR_unguarded(5) <= array_obj_ref_150_index_0_scale_req_1;
      reqR_unguarded(4) <= array_obj_ref_162_index_0_scale_req_1;
      reqR_unguarded(3) <= array_obj_ref_185_index_0_scale_req_1;
      reqR_unguarded(2) <= array_obj_ref_197_index_0_scale_req_1;
      reqR_unguarded(1) <= array_obj_ref_207_index_0_scale_req_1;
      reqR_unguarded(0) <= array_obj_ref_177_index_0_scale_req_1;
      array_obj_ref_125_index_0_scale_ack_1 <= ackR_unguarded(7);
      array_obj_ref_137_index_0_scale_ack_1 <= ackR_unguarded(6);
      array_obj_ref_150_index_0_scale_ack_1 <= ackR_unguarded(5);
      array_obj_ref_162_index_0_scale_ack_1 <= ackR_unguarded(4);
      array_obj_ref_185_index_0_scale_ack_1 <= ackR_unguarded(3);
      array_obj_ref_197_index_0_scale_ack_1 <= ackR_unguarded(2);
      array_obj_ref_207_index_0_scale_ack_1 <= ackR_unguarded(1);
      array_obj_ref_177_index_0_scale_ack_1 <= ackR_unguarded(0);
      ApIntMul_group_25_accessRegulator_0: access_regulator_base generic map (name => "ApIntMul_group_25_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      ApIntMul_group_25_accessRegulator_1: access_regulator_base generic map (name => "ApIntMul_group_25_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      ApIntMul_group_25_accessRegulator_2: access_regulator_base generic map (name => "ApIntMul_group_25_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      ApIntMul_group_25_accessRegulator_3: access_regulator_base generic map (name => "ApIntMul_group_25_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      ApIntMul_group_25_accessRegulator_4: access_regulator_base generic map (name => "ApIntMul_group_25_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      ApIntMul_group_25_accessRegulator_5: access_regulator_base generic map (name => "ApIntMul_group_25_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      ApIntMul_group_25_accessRegulator_6: access_regulator_base generic map (name => "ApIntMul_group_25_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      ApIntMul_group_25_accessRegulator_7: access_regulator_base generic map (name => "ApIntMul_group_25_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      ApIntMul_group_25_gI: SplitGuardInterface generic map(name => "ApIntMul_group_25_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          name => "ApIntMul_group_25",
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0100",
          constant_width => 4,
          use_constant  => true,
          full_rate  => false,
          no_arbitration => false,
          min_clock_period => false,
          num_reqs => 8,
          use_input_buffering => true,
          detailed_buffering_per_input => inBUFs,
          detailed_buffering_per_output => outBUFs --
        )
        port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : array_obj_ref_125_index_sum_1 
    ApIntAdd_group_26: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_output_port_124_scaled & R_input_port_123_scaled;
      array_obj_ref_125_index_partial_sum_1 <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_125_index_sum_1_req_0;
      array_obj_ref_125_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_125_index_sum_1_req_1;
      array_obj_ref_125_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_26_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_26_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_26",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 4, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : array_obj_ref_137_index_sum_1 
    ApIntAdd_group_27: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_output_port_136_scaled & R_input_port_135_scaled;
      array_obj_ref_137_index_partial_sum_1 <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_137_index_sum_1_req_0;
      array_obj_ref_137_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_137_index_sum_1_req_1;
      array_obj_ref_137_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_27_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_27_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_27",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 4, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : array_obj_ref_150_index_sum_1 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_output_port_149_scaled & R_input_port_148_scaled;
      array_obj_ref_150_index_partial_sum_1 <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_150_index_sum_1_req_0;
      array_obj_ref_150_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_150_index_sum_1_req_1;
      array_obj_ref_150_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 4, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_162_index_sum_1 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_output_port_161_scaled & R_input_port_160_scaled;
      array_obj_ref_162_index_partial_sum_1 <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_162_index_sum_1_req_0;
      array_obj_ref_162_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_162_index_sum_1_req_1;
      array_obj_ref_162_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 4, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : array_obj_ref_177_index_sum_1 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_output_port_176_scaled & R_input_port_175_scaled;
      array_obj_ref_177_index_partial_sum_1 <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_177_index_sum_1_req_0;
      array_obj_ref_177_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_177_index_sum_1_req_1;
      array_obj_ref_177_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 4, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : array_obj_ref_185_index_sum_1 
    ApIntAdd_group_31: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_output_port_184_scaled & R_input_port_183_scaled;
      array_obj_ref_185_index_partial_sum_1 <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_185_index_sum_1_req_0;
      array_obj_ref_185_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_185_index_sum_1_req_1;
      array_obj_ref_185_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_31_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_31_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 4, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : array_obj_ref_197_index_sum_1 
    ApIntAdd_group_32: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_output_port_196_scaled & R_input_port_195_scaled;
      array_obj_ref_197_index_partial_sum_1 <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_197_index_sum_1_req_0;
      array_obj_ref_197_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_197_index_sum_1_req_1;
      array_obj_ref_197_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_32_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_32_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_32",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 4, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared split operator group (33) : array_obj_ref_207_index_sum_1 
    ApIntAdd_group_33: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_output_port_206_scaled & R_input_port_205_scaled;
      array_obj_ref_207_index_partial_sum_1 <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_207_index_sum_1_req_0;
      array_obj_ref_207_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_207_index_sum_1_req_1;
      array_obj_ref_207_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_33_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_33_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_33",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 4, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared load operator group (0) : array_obj_ref_125_load_0 array_obj_ref_137_load_0 array_obj_ref_150_load_0 array_obj_ref_162_load_0 array_obj_ref_185_load_0 array_obj_ref_197_load_0 array_obj_ref_207_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 6 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 6 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant inBUFs : IntegerArray(6 downto 0) := (6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(6 downto 0) := (6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      reqL_unguarded(6) <= array_obj_ref_125_load_0_req_0;
      reqL_unguarded(5) <= array_obj_ref_137_load_0_req_0;
      reqL_unguarded(4) <= array_obj_ref_150_load_0_req_0;
      reqL_unguarded(3) <= array_obj_ref_162_load_0_req_0;
      reqL_unguarded(2) <= array_obj_ref_185_load_0_req_0;
      reqL_unguarded(1) <= array_obj_ref_197_load_0_req_0;
      reqL_unguarded(0) <= array_obj_ref_207_load_0_req_0;
      array_obj_ref_125_load_0_ack_0 <= ackL_unguarded(6);
      array_obj_ref_137_load_0_ack_0 <= ackL_unguarded(5);
      array_obj_ref_150_load_0_ack_0 <= ackL_unguarded(4);
      array_obj_ref_162_load_0_ack_0 <= ackL_unguarded(3);
      array_obj_ref_185_load_0_ack_0 <= ackL_unguarded(2);
      array_obj_ref_197_load_0_ack_0 <= ackL_unguarded(1);
      array_obj_ref_207_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(6) <= array_obj_ref_125_load_0_req_1;
      reqR_unguarded(5) <= array_obj_ref_137_load_0_req_1;
      reqR_unguarded(4) <= array_obj_ref_150_load_0_req_1;
      reqR_unguarded(3) <= array_obj_ref_162_load_0_req_1;
      reqR_unguarded(2) <= array_obj_ref_185_load_0_req_1;
      reqR_unguarded(1) <= array_obj_ref_197_load_0_req_1;
      reqR_unguarded(0) <= array_obj_ref_207_load_0_req_1;
      array_obj_ref_125_load_0_ack_1 <= ackR_unguarded(6);
      array_obj_ref_137_load_0_ack_1 <= ackR_unguarded(5);
      array_obj_ref_150_load_0_ack_1 <= ackR_unguarded(4);
      array_obj_ref_162_load_0_ack_1 <= ackR_unguarded(3);
      array_obj_ref_185_load_0_ack_1 <= ackR_unguarded(2);
      array_obj_ref_197_load_0_ack_1 <= ackR_unguarded(1);
      array_obj_ref_207_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_125_word_address_0 & array_obj_ref_137_word_address_0 & array_obj_ref_150_word_address_0 & array_obj_ref_162_word_address_0 & array_obj_ref_185_word_address_0 & array_obj_ref_197_word_address_0 & array_obj_ref_207_word_address_0;
      array_obj_ref_125_data_0 <= data_out(13 downto 12);
      array_obj_ref_137_data_0 <= data_out(11 downto 10);
      array_obj_ref_150_data_0 <= data_out(9 downto 8);
      array_obj_ref_162_data_0 <= data_out(7 downto 6);
      array_obj_ref_185_data_0 <= data_out(5 downto 4);
      array_obj_ref_197_data_0 <= data_out(3 downto 2);
      array_obj_ref_207_data_0 <= data_out(1 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 4,
        num_reqs => 7,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(3 downto 0),
          mtag => memory_space_0_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 2,
        num_reqs => 7,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(1 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : array_obj_ref_177_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(3 downto 0);
      signal data_in: std_logic_vector(1 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_177_store_0_req_0;
      array_obj_ref_177_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_177_store_0_req_1;
      array_obj_ref_177_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_177_word_address_0;
      data_in <= array_obj_ref_177_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 4,
        data_width => 2,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(3 downto 0),
          mdata => memory_space_0_sr_data(1 downto 0),
          mtag => memory_space_0_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end updateCounter_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    initialiseCounters_tag_in: in std_logic_vector(1 downto 0);
    initialiseCounters_tag_out: out std_logic_vector(1 downto 0);
    initialiseCounters_start_req : in std_logic;
    initialiseCounters_start_ack : out std_logic;
    initialiseCounters_fin_req   : in std_logic;
    initialiseCounters_fin_ack   : out std_logic;
    clk : in std_logic;
    reset : in std_logic;
    in_data_1_pipe_write_data: in std_logic_vector(31 downto 0);
    in_data_1_pipe_write_req : in std_logic_vector(0 downto 0);
    in_data_1_pipe_write_ack : out std_logic_vector(0 downto 0);
    in_data_2_pipe_write_data: in std_logic_vector(31 downto 0);
    in_data_2_pipe_write_req : in std_logic_vector(0 downto 0);
    in_data_2_pipe_write_ack : out std_logic_vector(0 downto 0);
    in_data_3_pipe_write_data: in std_logic_vector(31 downto 0);
    in_data_3_pipe_write_req : in std_logic_vector(0 downto 0);
    in_data_3_pipe_write_ack : out std_logic_vector(0 downto 0);
    in_data_4_pipe_write_data: in std_logic_vector(31 downto 0);
    in_data_4_pipe_write_req : in std_logic_vector(0 downto 0);
    in_data_4_pipe_write_ack : out std_logic_vector(0 downto 0);
    out_data_1_pipe_read_data: out std_logic_vector(31 downto 0);
    out_data_1_pipe_read_req : in std_logic_vector(0 downto 0);
    out_data_1_pipe_read_ack : out std_logic_vector(0 downto 0);
    out_data_2_pipe_read_data: out std_logic_vector(31 downto 0);
    out_data_2_pipe_read_req : in std_logic_vector(0 downto 0);
    out_data_2_pipe_read_ack : out std_logic_vector(0 downto 0);
    out_data_3_pipe_read_data: out std_logic_vector(31 downto 0);
    out_data_3_pipe_read_req : in std_logic_vector(0 downto 0);
    out_data_3_pipe_read_ack : out std_logic_vector(0 downto 0);
    out_data_4_pipe_read_data: out std_logic_vector(31 downto 0);
    out_data_4_pipe_read_req : in std_logic_vector(0 downto 0);
    out_data_4_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(3 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(19 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(1 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(1 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(1 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(7 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(3 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(39 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(1 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(5 downto 0);
  -- declarations related to module initialiseCounters
  component initialiseCounters is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(1 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- declarations related to module inputPort_1_Daemon
  component inputPort_1_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      in_data_1_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_1_pipe_read_data : in   std_logic_vector(31 downto 0);
      noblock_obuf_1_3_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_3_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_1_4_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_4_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_1_1_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_1_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_1_2_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_2_pipe_write_data : out  std_logic_vector(32 downto 0);
      updateCounter_call_reqs : out  std_logic_vector(0 downto 0);
      updateCounter_call_acks : in   std_logic_vector(0 downto 0);
      updateCounter_call_data : out  std_logic_vector(16 downto 0);
      updateCounter_call_tag  :  out  std_logic_vector(0 downto 0);
      updateCounter_return_reqs : out  std_logic_vector(0 downto 0);
      updateCounter_return_acks : in   std_logic_vector(0 downto 0);
      updateCounter_return_data : in   std_logic_vector(0 downto 0);
      updateCounter_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module inputPort_1_Daemon
  signal inputPort_1_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal inputPort_1_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal inputPort_1_Daemon_start_req : std_logic;
  signal inputPort_1_Daemon_start_ack : std_logic;
  signal inputPort_1_Daemon_fin_req   : std_logic;
  signal inputPort_1_Daemon_fin_ack : std_logic;
  -- declarations related to module inputPort_2_Daemon
  component inputPort_2_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      in_data_2_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_2_pipe_read_data : in   std_logic_vector(31 downto 0);
      noblock_obuf_2_1_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_1_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_2_2_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_2_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_2_3_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_3_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_2_4_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_4_pipe_write_data : out  std_logic_vector(32 downto 0);
      updateCounter_call_reqs : out  std_logic_vector(0 downto 0);
      updateCounter_call_acks : in   std_logic_vector(0 downto 0);
      updateCounter_call_data : out  std_logic_vector(16 downto 0);
      updateCounter_call_tag  :  out  std_logic_vector(0 downto 0);
      updateCounter_return_reqs : out  std_logic_vector(0 downto 0);
      updateCounter_return_acks : in   std_logic_vector(0 downto 0);
      updateCounter_return_data : in   std_logic_vector(0 downto 0);
      updateCounter_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module inputPort_2_Daemon
  signal inputPort_2_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal inputPort_2_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal inputPort_2_Daemon_start_req : std_logic;
  signal inputPort_2_Daemon_start_ack : std_logic;
  signal inputPort_2_Daemon_fin_req   : std_logic;
  signal inputPort_2_Daemon_fin_ack : std_logic;
  -- declarations related to module inputPort_3_Daemon
  component inputPort_3_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      in_data_3_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_3_pipe_read_data : in   std_logic_vector(31 downto 0);
      noblock_obuf_3_2_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_2_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_3_3_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_3_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_3_4_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_4_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_3_1_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_1_pipe_write_data : out  std_logic_vector(32 downto 0);
      updateCounter_call_reqs : out  std_logic_vector(0 downto 0);
      updateCounter_call_acks : in   std_logic_vector(0 downto 0);
      updateCounter_call_data : out  std_logic_vector(16 downto 0);
      updateCounter_call_tag  :  out  std_logic_vector(0 downto 0);
      updateCounter_return_reqs : out  std_logic_vector(0 downto 0);
      updateCounter_return_acks : in   std_logic_vector(0 downto 0);
      updateCounter_return_data : in   std_logic_vector(0 downto 0);
      updateCounter_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module inputPort_3_Daemon
  signal inputPort_3_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal inputPort_3_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal inputPort_3_Daemon_start_req : std_logic;
  signal inputPort_3_Daemon_start_ack : std_logic;
  signal inputPort_3_Daemon_fin_req   : std_logic;
  signal inputPort_3_Daemon_fin_ack : std_logic;
  -- declarations related to module inputPort_4_Daemon
  component inputPort_4_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      in_data_4_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_4_pipe_read_data : in   std_logic_vector(31 downto 0);
      noblock_obuf_4_1_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_1_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_4_2_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_2_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_4_3_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_3_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_4_4_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_4_pipe_write_data : out  std_logic_vector(32 downto 0);
      updateCounter_call_reqs : out  std_logic_vector(0 downto 0);
      updateCounter_call_acks : in   std_logic_vector(0 downto 0);
      updateCounter_call_data : out  std_logic_vector(16 downto 0);
      updateCounter_call_tag  :  out  std_logic_vector(0 downto 0);
      updateCounter_return_reqs : out  std_logic_vector(0 downto 0);
      updateCounter_return_acks : in   std_logic_vector(0 downto 0);
      updateCounter_return_data : in   std_logic_vector(0 downto 0);
      updateCounter_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module inputPort_4_Daemon
  signal inputPort_4_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal inputPort_4_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal inputPort_4_Daemon_start_req : std_logic;
  signal inputPort_4_Daemon_start_ack : std_logic;
  signal inputPort_4_Daemon_fin_req   : std_logic;
  signal inputPort_4_Daemon_fin_ack : std_logic;
  -- declarations related to module outputPort_1_Daemon
  component outputPort_1_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      noblock_obuf_4_1_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_1_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_2_1_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_1_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_1_1_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_1_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_3_1_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_1_pipe_read_data : in   std_logic_vector(32 downto 0);
      out_data_1_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_data_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_data_1_pipe_write_data : out  std_logic_vector(31 downto 0);
      updateCounter_call_reqs : out  std_logic_vector(0 downto 0);
      updateCounter_call_acks : in   std_logic_vector(0 downto 0);
      updateCounter_call_data : out  std_logic_vector(16 downto 0);
      updateCounter_call_tag  :  out  std_logic_vector(0 downto 0);
      updateCounter_return_reqs : out  std_logic_vector(0 downto 0);
      updateCounter_return_acks : in   std_logic_vector(0 downto 0);
      updateCounter_return_data : in   std_logic_vector(0 downto 0);
      updateCounter_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module outputPort_1_Daemon
  signal outputPort_1_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal outputPort_1_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal outputPort_1_Daemon_start_req : std_logic;
  signal outputPort_1_Daemon_start_ack : std_logic;
  signal outputPort_1_Daemon_fin_req   : std_logic;
  signal outputPort_1_Daemon_fin_ack : std_logic;
  -- declarations related to module outputPort_2_Daemon
  component outputPort_2_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      noblock_obuf_1_2_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_2_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_3_2_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_2_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_4_2_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_2_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_2_2_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_2_pipe_read_data : in   std_logic_vector(32 downto 0);
      out_data_2_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_data_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_data_2_pipe_write_data : out  std_logic_vector(31 downto 0);
      updateCounter_call_reqs : out  std_logic_vector(0 downto 0);
      updateCounter_call_acks : in   std_logic_vector(0 downto 0);
      updateCounter_call_data : out  std_logic_vector(16 downto 0);
      updateCounter_call_tag  :  out  std_logic_vector(0 downto 0);
      updateCounter_return_reqs : out  std_logic_vector(0 downto 0);
      updateCounter_return_acks : in   std_logic_vector(0 downto 0);
      updateCounter_return_data : in   std_logic_vector(0 downto 0);
      updateCounter_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module outputPort_2_Daemon
  signal outputPort_2_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal outputPort_2_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal outputPort_2_Daemon_start_req : std_logic;
  signal outputPort_2_Daemon_start_ack : std_logic;
  signal outputPort_2_Daemon_fin_req   : std_logic;
  signal outputPort_2_Daemon_fin_ack : std_logic;
  -- declarations related to module outputPort_3_Daemon
  component outputPort_3_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      noblock_obuf_1_3_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_3_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_3_3_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_3_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_4_3_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_3_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_2_3_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_3_pipe_read_data : in   std_logic_vector(32 downto 0);
      out_data_3_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_data_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_data_3_pipe_write_data : out  std_logic_vector(31 downto 0);
      updateCounter_call_reqs : out  std_logic_vector(0 downto 0);
      updateCounter_call_acks : in   std_logic_vector(0 downto 0);
      updateCounter_call_data : out  std_logic_vector(16 downto 0);
      updateCounter_call_tag  :  out  std_logic_vector(0 downto 0);
      updateCounter_return_reqs : out  std_logic_vector(0 downto 0);
      updateCounter_return_acks : in   std_logic_vector(0 downto 0);
      updateCounter_return_data : in   std_logic_vector(0 downto 0);
      updateCounter_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module outputPort_3_Daemon
  signal outputPort_3_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal outputPort_3_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal outputPort_3_Daemon_start_req : std_logic;
  signal outputPort_3_Daemon_start_ack : std_logic;
  signal outputPort_3_Daemon_fin_req   : std_logic;
  signal outputPort_3_Daemon_fin_ack : std_logic;
  -- declarations related to module outputPort_4_Daemon
  component outputPort_4_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      noblock_obuf_1_4_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_4_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_3_4_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_4_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_2_4_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_4_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_4_4_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_4_pipe_read_data : in   std_logic_vector(32 downto 0);
      out_data_4_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_data_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_data_4_pipe_write_data : out  std_logic_vector(31 downto 0);
      updateCounter_call_reqs : out  std_logic_vector(0 downto 0);
      updateCounter_call_acks : in   std_logic_vector(0 downto 0);
      updateCounter_call_data : out  std_logic_vector(16 downto 0);
      updateCounter_call_tag  :  out  std_logic_vector(0 downto 0);
      updateCounter_return_reqs : out  std_logic_vector(0 downto 0);
      updateCounter_return_acks : in   std_logic_vector(0 downto 0);
      updateCounter_return_data : in   std_logic_vector(0 downto 0);
      updateCounter_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module outputPort_4_Daemon
  signal outputPort_4_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal outputPort_4_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal outputPort_4_Daemon_start_req : std_logic;
  signal outputPort_4_Daemon_start_ack : std_logic;
  signal outputPort_4_Daemon_fin_req   : std_logic;
  signal outputPort_4_Daemon_fin_ack : std_logic;
  -- declarations related to module prioritySelect
  -- declarations related to module updateCounter
  component updateCounter is -- 
    generic (tag_length : integer); 
    port ( -- 
      input_port : in  std_logic_vector(7 downto 0);
      output_port : in  std_logic_vector(7 downto 0);
      up : in  std_logic_vector(0 downto 0);
      continue : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(3 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(1 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(1 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module updateCounter
  signal updateCounter_input_port :  std_logic_vector(7 downto 0);
  signal updateCounter_output_port :  std_logic_vector(7 downto 0);
  signal updateCounter_up :  std_logic_vector(0 downto 0);
  signal updateCounter_continue :  std_logic_vector(0 downto 0);
  signal updateCounter_in_args    : std_logic_vector(16 downto 0);
  signal updateCounter_out_args   : std_logic_vector(0 downto 0);
  signal updateCounter_tag_in    : std_logic_vector(4 downto 0) := (others => '0');
  signal updateCounter_tag_out   : std_logic_vector(4 downto 0);
  signal updateCounter_start_req : std_logic;
  signal updateCounter_start_ack : std_logic;
  signal updateCounter_fin_req   : std_logic;
  signal updateCounter_fin_ack : std_logic;
  -- caller side aggregated signals for module updateCounter
  signal updateCounter_call_reqs: std_logic_vector(7 downto 0);
  signal updateCounter_call_acks: std_logic_vector(7 downto 0);
  signal updateCounter_return_reqs: std_logic_vector(7 downto 0);
  signal updateCounter_return_acks: std_logic_vector(7 downto 0);
  signal updateCounter_call_data: std_logic_vector(135 downto 0);
  signal updateCounter_call_tag: std_logic_vector(7 downto 0);
  signal updateCounter_return_data: std_logic_vector(7 downto 0);
  signal updateCounter_return_tag: std_logic_vector(7 downto 0);
  -- aggregate signals for read from pipe in_data_1
  signal in_data_1_pipe_read_data: std_logic_vector(31 downto 0);
  signal in_data_1_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_data_1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe in_data_2
  signal in_data_2_pipe_read_data: std_logic_vector(31 downto 0);
  signal in_data_2_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_data_2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe in_data_3
  signal in_data_3_pipe_read_data: std_logic_vector(31 downto 0);
  signal in_data_3_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_data_3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe in_data_4
  signal in_data_4_pipe_read_data: std_logic_vector(31 downto 0);
  signal in_data_4_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_data_4_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_1_1
  signal noblock_obuf_1_1_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_1_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_1_1
  signal noblock_obuf_1_1_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_1_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_1_2
  signal noblock_obuf_1_2_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_2_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_1_2
  signal noblock_obuf_1_2_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_2_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_1_3
  signal noblock_obuf_1_3_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_3_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_1_3
  signal noblock_obuf_1_3_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_3_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_1_4
  signal noblock_obuf_1_4_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_4_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_4_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_1_4
  signal noblock_obuf_1_4_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_4_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_4_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_2_1
  signal noblock_obuf_2_1_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_1_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_2_1
  signal noblock_obuf_2_1_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_1_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_2_2
  signal noblock_obuf_2_2_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_2_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_2_2
  signal noblock_obuf_2_2_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_2_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_2_3
  signal noblock_obuf_2_3_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_3_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_2_3
  signal noblock_obuf_2_3_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_3_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_2_4
  signal noblock_obuf_2_4_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_4_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_4_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_2_4
  signal noblock_obuf_2_4_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_4_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_4_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_3_1
  signal noblock_obuf_3_1_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_1_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_3_1
  signal noblock_obuf_3_1_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_1_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_3_2
  signal noblock_obuf_3_2_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_2_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_3_2
  signal noblock_obuf_3_2_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_2_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_3_3
  signal noblock_obuf_3_3_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_3_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_3_3
  signal noblock_obuf_3_3_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_3_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_3_4
  signal noblock_obuf_3_4_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_4_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_4_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_3_4
  signal noblock_obuf_3_4_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_4_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_4_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_4_1
  signal noblock_obuf_4_1_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_1_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_4_1
  signal noblock_obuf_4_1_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_1_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_4_2
  signal noblock_obuf_4_2_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_2_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_4_2
  signal noblock_obuf_4_2_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_2_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_4_3
  signal noblock_obuf_4_3_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_3_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_4_3
  signal noblock_obuf_4_3_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_3_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_4_4
  signal noblock_obuf_4_4_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_4_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_4_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_4_4
  signal noblock_obuf_4_4_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_4_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_4_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_data_1
  signal out_data_1_pipe_write_data: std_logic_vector(31 downto 0);
  signal out_data_1_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_data_1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_data_2
  signal out_data_2_pipe_write_data: std_logic_vector(31 downto 0);
  signal out_data_2_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_data_2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_data_3
  signal out_data_3_pipe_write_data: std_logic_vector(31 downto 0);
  signal out_data_3_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_data_3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_data_4
  signal out_data_4_pipe_write_data: std_logic_vector(31 downto 0);
  signal out_data_4_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_data_4_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module initialiseCounters
  initialiseCounters_instance:initialiseCounters-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => initialiseCounters_start_req,
      start_ack => initialiseCounters_start_ack,
      fin_req => initialiseCounters_fin_req,
      fin_ack => initialiseCounters_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_sr_req => memory_space_0_sr_req(1 downto 1),
      memory_space_0_sr_ack => memory_space_0_sr_ack(1 downto 1),
      memory_space_0_sr_addr => memory_space_0_sr_addr(7 downto 4),
      memory_space_0_sr_data => memory_space_0_sr_data(3 downto 2),
      memory_space_0_sr_tag => memory_space_0_sr_tag(39 downto 20),
      memory_space_0_sc_req => memory_space_0_sc_req(1 downto 1),
      memory_space_0_sc_ack => memory_space_0_sc_ack(1 downto 1),
      memory_space_0_sc_tag => memory_space_0_sc_tag(5 downto 3),
      tag_in => initialiseCounters_tag_in,
      tag_out => initialiseCounters_tag_out-- 
    ); -- 
  -- module inputPort_1_Daemon
  inputPort_1_Daemon_instance:inputPort_1_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => inputPort_1_Daemon_start_req,
      start_ack => inputPort_1_Daemon_start_ack,
      fin_req => inputPort_1_Daemon_fin_req,
      fin_ack => inputPort_1_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      in_data_1_pipe_read_req => in_data_1_pipe_read_req(0 downto 0),
      in_data_1_pipe_read_ack => in_data_1_pipe_read_ack(0 downto 0),
      in_data_1_pipe_read_data => in_data_1_pipe_read_data(31 downto 0),
      noblock_obuf_1_3_pipe_write_req => noblock_obuf_1_3_pipe_write_req(0 downto 0),
      noblock_obuf_1_3_pipe_write_ack => noblock_obuf_1_3_pipe_write_ack(0 downto 0),
      noblock_obuf_1_3_pipe_write_data => noblock_obuf_1_3_pipe_write_data(32 downto 0),
      noblock_obuf_1_4_pipe_write_req => noblock_obuf_1_4_pipe_write_req(0 downto 0),
      noblock_obuf_1_4_pipe_write_ack => noblock_obuf_1_4_pipe_write_ack(0 downto 0),
      noblock_obuf_1_4_pipe_write_data => noblock_obuf_1_4_pipe_write_data(32 downto 0),
      noblock_obuf_1_1_pipe_write_req => noblock_obuf_1_1_pipe_write_req(0 downto 0),
      noblock_obuf_1_1_pipe_write_ack => noblock_obuf_1_1_pipe_write_ack(0 downto 0),
      noblock_obuf_1_1_pipe_write_data => noblock_obuf_1_1_pipe_write_data(32 downto 0),
      noblock_obuf_1_2_pipe_write_req => noblock_obuf_1_2_pipe_write_req(0 downto 0),
      noblock_obuf_1_2_pipe_write_ack => noblock_obuf_1_2_pipe_write_ack(0 downto 0),
      noblock_obuf_1_2_pipe_write_data => noblock_obuf_1_2_pipe_write_data(32 downto 0),
      updateCounter_call_reqs => updateCounter_call_reqs(7 downto 7),
      updateCounter_call_acks => updateCounter_call_acks(7 downto 7),
      updateCounter_call_data => updateCounter_call_data(135 downto 119),
      updateCounter_call_tag => updateCounter_call_tag(7 downto 7),
      updateCounter_return_reqs => updateCounter_return_reqs(7 downto 7),
      updateCounter_return_acks => updateCounter_return_acks(7 downto 7),
      updateCounter_return_data => updateCounter_return_data(7 downto 7),
      updateCounter_return_tag => updateCounter_return_tag(7 downto 7),
      tag_in => inputPort_1_Daemon_tag_in,
      tag_out => inputPort_1_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  inputPort_1_Daemon_tag_in <= (others => '0');
  inputPort_1_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => inputPort_1_Daemon_start_req, start_ack => inputPort_1_Daemon_start_ack,  fin_req => inputPort_1_Daemon_fin_req,  fin_ack => inputPort_1_Daemon_fin_ack);
  -- module inputPort_2_Daemon
  inputPort_2_Daemon_instance:inputPort_2_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => inputPort_2_Daemon_start_req,
      start_ack => inputPort_2_Daemon_start_ack,
      fin_req => inputPort_2_Daemon_fin_req,
      fin_ack => inputPort_2_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      in_data_2_pipe_read_req => in_data_2_pipe_read_req(0 downto 0),
      in_data_2_pipe_read_ack => in_data_2_pipe_read_ack(0 downto 0),
      in_data_2_pipe_read_data => in_data_2_pipe_read_data(31 downto 0),
      noblock_obuf_2_1_pipe_write_req => noblock_obuf_2_1_pipe_write_req(0 downto 0),
      noblock_obuf_2_1_pipe_write_ack => noblock_obuf_2_1_pipe_write_ack(0 downto 0),
      noblock_obuf_2_1_pipe_write_data => noblock_obuf_2_1_pipe_write_data(32 downto 0),
      noblock_obuf_2_2_pipe_write_req => noblock_obuf_2_2_pipe_write_req(0 downto 0),
      noblock_obuf_2_2_pipe_write_ack => noblock_obuf_2_2_pipe_write_ack(0 downto 0),
      noblock_obuf_2_2_pipe_write_data => noblock_obuf_2_2_pipe_write_data(32 downto 0),
      noblock_obuf_2_3_pipe_write_req => noblock_obuf_2_3_pipe_write_req(0 downto 0),
      noblock_obuf_2_3_pipe_write_ack => noblock_obuf_2_3_pipe_write_ack(0 downto 0),
      noblock_obuf_2_3_pipe_write_data => noblock_obuf_2_3_pipe_write_data(32 downto 0),
      noblock_obuf_2_4_pipe_write_req => noblock_obuf_2_4_pipe_write_req(0 downto 0),
      noblock_obuf_2_4_pipe_write_ack => noblock_obuf_2_4_pipe_write_ack(0 downto 0),
      noblock_obuf_2_4_pipe_write_data => noblock_obuf_2_4_pipe_write_data(32 downto 0),
      updateCounter_call_reqs => updateCounter_call_reqs(6 downto 6),
      updateCounter_call_acks => updateCounter_call_acks(6 downto 6),
      updateCounter_call_data => updateCounter_call_data(118 downto 102),
      updateCounter_call_tag => updateCounter_call_tag(6 downto 6),
      updateCounter_return_reqs => updateCounter_return_reqs(6 downto 6),
      updateCounter_return_acks => updateCounter_return_acks(6 downto 6),
      updateCounter_return_data => updateCounter_return_data(6 downto 6),
      updateCounter_return_tag => updateCounter_return_tag(6 downto 6),
      tag_in => inputPort_2_Daemon_tag_in,
      tag_out => inputPort_2_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  inputPort_2_Daemon_tag_in <= (others => '0');
  inputPort_2_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => inputPort_2_Daemon_start_req, start_ack => inputPort_2_Daemon_start_ack,  fin_req => inputPort_2_Daemon_fin_req,  fin_ack => inputPort_2_Daemon_fin_ack);
  -- module inputPort_3_Daemon
  inputPort_3_Daemon_instance:inputPort_3_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => inputPort_3_Daemon_start_req,
      start_ack => inputPort_3_Daemon_start_ack,
      fin_req => inputPort_3_Daemon_fin_req,
      fin_ack => inputPort_3_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      in_data_3_pipe_read_req => in_data_3_pipe_read_req(0 downto 0),
      in_data_3_pipe_read_ack => in_data_3_pipe_read_ack(0 downto 0),
      in_data_3_pipe_read_data => in_data_3_pipe_read_data(31 downto 0),
      noblock_obuf_3_2_pipe_write_req => noblock_obuf_3_2_pipe_write_req(0 downto 0),
      noblock_obuf_3_2_pipe_write_ack => noblock_obuf_3_2_pipe_write_ack(0 downto 0),
      noblock_obuf_3_2_pipe_write_data => noblock_obuf_3_2_pipe_write_data(32 downto 0),
      noblock_obuf_3_3_pipe_write_req => noblock_obuf_3_3_pipe_write_req(0 downto 0),
      noblock_obuf_3_3_pipe_write_ack => noblock_obuf_3_3_pipe_write_ack(0 downto 0),
      noblock_obuf_3_3_pipe_write_data => noblock_obuf_3_3_pipe_write_data(32 downto 0),
      noblock_obuf_3_4_pipe_write_req => noblock_obuf_3_4_pipe_write_req(0 downto 0),
      noblock_obuf_3_4_pipe_write_ack => noblock_obuf_3_4_pipe_write_ack(0 downto 0),
      noblock_obuf_3_4_pipe_write_data => noblock_obuf_3_4_pipe_write_data(32 downto 0),
      noblock_obuf_3_1_pipe_write_req => noblock_obuf_3_1_pipe_write_req(0 downto 0),
      noblock_obuf_3_1_pipe_write_ack => noblock_obuf_3_1_pipe_write_ack(0 downto 0),
      noblock_obuf_3_1_pipe_write_data => noblock_obuf_3_1_pipe_write_data(32 downto 0),
      updateCounter_call_reqs => updateCounter_call_reqs(5 downto 5),
      updateCounter_call_acks => updateCounter_call_acks(5 downto 5),
      updateCounter_call_data => updateCounter_call_data(101 downto 85),
      updateCounter_call_tag => updateCounter_call_tag(5 downto 5),
      updateCounter_return_reqs => updateCounter_return_reqs(5 downto 5),
      updateCounter_return_acks => updateCounter_return_acks(5 downto 5),
      updateCounter_return_data => updateCounter_return_data(5 downto 5),
      updateCounter_return_tag => updateCounter_return_tag(5 downto 5),
      tag_in => inputPort_3_Daemon_tag_in,
      tag_out => inputPort_3_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  inputPort_3_Daemon_tag_in <= (others => '0');
  inputPort_3_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => inputPort_3_Daemon_start_req, start_ack => inputPort_3_Daemon_start_ack,  fin_req => inputPort_3_Daemon_fin_req,  fin_ack => inputPort_3_Daemon_fin_ack);
  -- module inputPort_4_Daemon
  inputPort_4_Daemon_instance:inputPort_4_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => inputPort_4_Daemon_start_req,
      start_ack => inputPort_4_Daemon_start_ack,
      fin_req => inputPort_4_Daemon_fin_req,
      fin_ack => inputPort_4_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      in_data_4_pipe_read_req => in_data_4_pipe_read_req(0 downto 0),
      in_data_4_pipe_read_ack => in_data_4_pipe_read_ack(0 downto 0),
      in_data_4_pipe_read_data => in_data_4_pipe_read_data(31 downto 0),
      noblock_obuf_4_1_pipe_write_req => noblock_obuf_4_1_pipe_write_req(0 downto 0),
      noblock_obuf_4_1_pipe_write_ack => noblock_obuf_4_1_pipe_write_ack(0 downto 0),
      noblock_obuf_4_1_pipe_write_data => noblock_obuf_4_1_pipe_write_data(32 downto 0),
      noblock_obuf_4_2_pipe_write_req => noblock_obuf_4_2_pipe_write_req(0 downto 0),
      noblock_obuf_4_2_pipe_write_ack => noblock_obuf_4_2_pipe_write_ack(0 downto 0),
      noblock_obuf_4_2_pipe_write_data => noblock_obuf_4_2_pipe_write_data(32 downto 0),
      noblock_obuf_4_3_pipe_write_req => noblock_obuf_4_3_pipe_write_req(0 downto 0),
      noblock_obuf_4_3_pipe_write_ack => noblock_obuf_4_3_pipe_write_ack(0 downto 0),
      noblock_obuf_4_3_pipe_write_data => noblock_obuf_4_3_pipe_write_data(32 downto 0),
      noblock_obuf_4_4_pipe_write_req => noblock_obuf_4_4_pipe_write_req(0 downto 0),
      noblock_obuf_4_4_pipe_write_ack => noblock_obuf_4_4_pipe_write_ack(0 downto 0),
      noblock_obuf_4_4_pipe_write_data => noblock_obuf_4_4_pipe_write_data(32 downto 0),
      updateCounter_call_reqs => updateCounter_call_reqs(4 downto 4),
      updateCounter_call_acks => updateCounter_call_acks(4 downto 4),
      updateCounter_call_data => updateCounter_call_data(84 downto 68),
      updateCounter_call_tag => updateCounter_call_tag(4 downto 4),
      updateCounter_return_reqs => updateCounter_return_reqs(4 downto 4),
      updateCounter_return_acks => updateCounter_return_acks(4 downto 4),
      updateCounter_return_data => updateCounter_return_data(4 downto 4),
      updateCounter_return_tag => updateCounter_return_tag(4 downto 4),
      tag_in => inputPort_4_Daemon_tag_in,
      tag_out => inputPort_4_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  inputPort_4_Daemon_tag_in <= (others => '0');
  inputPort_4_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => inputPort_4_Daemon_start_req, start_ack => inputPort_4_Daemon_start_ack,  fin_req => inputPort_4_Daemon_fin_req,  fin_ack => inputPort_4_Daemon_fin_ack);
  -- module outputPort_1_Daemon
  outputPort_1_Daemon_instance:outputPort_1_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => outputPort_1_Daemon_start_req,
      start_ack => outputPort_1_Daemon_start_ack,
      fin_req => outputPort_1_Daemon_fin_req,
      fin_ack => outputPort_1_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      noblock_obuf_4_1_pipe_read_req => noblock_obuf_4_1_pipe_read_req(0 downto 0),
      noblock_obuf_4_1_pipe_read_ack => noblock_obuf_4_1_pipe_read_ack(0 downto 0),
      noblock_obuf_4_1_pipe_read_data => noblock_obuf_4_1_pipe_read_data(32 downto 0),
      noblock_obuf_2_1_pipe_read_req => noblock_obuf_2_1_pipe_read_req(0 downto 0),
      noblock_obuf_2_1_pipe_read_ack => noblock_obuf_2_1_pipe_read_ack(0 downto 0),
      noblock_obuf_2_1_pipe_read_data => noblock_obuf_2_1_pipe_read_data(32 downto 0),
      noblock_obuf_1_1_pipe_read_req => noblock_obuf_1_1_pipe_read_req(0 downto 0),
      noblock_obuf_1_1_pipe_read_ack => noblock_obuf_1_1_pipe_read_ack(0 downto 0),
      noblock_obuf_1_1_pipe_read_data => noblock_obuf_1_1_pipe_read_data(32 downto 0),
      noblock_obuf_3_1_pipe_read_req => noblock_obuf_3_1_pipe_read_req(0 downto 0),
      noblock_obuf_3_1_pipe_read_ack => noblock_obuf_3_1_pipe_read_ack(0 downto 0),
      noblock_obuf_3_1_pipe_read_data => noblock_obuf_3_1_pipe_read_data(32 downto 0),
      out_data_1_pipe_write_req => out_data_1_pipe_write_req(0 downto 0),
      out_data_1_pipe_write_ack => out_data_1_pipe_write_ack(0 downto 0),
      out_data_1_pipe_write_data => out_data_1_pipe_write_data(31 downto 0),
      updateCounter_call_reqs => updateCounter_call_reqs(2 downto 2),
      updateCounter_call_acks => updateCounter_call_acks(2 downto 2),
      updateCounter_call_data => updateCounter_call_data(50 downto 34),
      updateCounter_call_tag => updateCounter_call_tag(2 downto 2),
      updateCounter_return_reqs => updateCounter_return_reqs(2 downto 2),
      updateCounter_return_acks => updateCounter_return_acks(2 downto 2),
      updateCounter_return_data => updateCounter_return_data(2 downto 2),
      updateCounter_return_tag => updateCounter_return_tag(2 downto 2),
      tag_in => outputPort_1_Daemon_tag_in,
      tag_out => outputPort_1_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  outputPort_1_Daemon_tag_in <= (others => '0');
  outputPort_1_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => outputPort_1_Daemon_start_req, start_ack => outputPort_1_Daemon_start_ack,  fin_req => outputPort_1_Daemon_fin_req,  fin_ack => outputPort_1_Daemon_fin_ack);
  -- module outputPort_2_Daemon
  outputPort_2_Daemon_instance:outputPort_2_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => outputPort_2_Daemon_start_req,
      start_ack => outputPort_2_Daemon_start_ack,
      fin_req => outputPort_2_Daemon_fin_req,
      fin_ack => outputPort_2_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      noblock_obuf_1_2_pipe_read_req => noblock_obuf_1_2_pipe_read_req(0 downto 0),
      noblock_obuf_1_2_pipe_read_ack => noblock_obuf_1_2_pipe_read_ack(0 downto 0),
      noblock_obuf_1_2_pipe_read_data => noblock_obuf_1_2_pipe_read_data(32 downto 0),
      noblock_obuf_3_2_pipe_read_req => noblock_obuf_3_2_pipe_read_req(0 downto 0),
      noblock_obuf_3_2_pipe_read_ack => noblock_obuf_3_2_pipe_read_ack(0 downto 0),
      noblock_obuf_3_2_pipe_read_data => noblock_obuf_3_2_pipe_read_data(32 downto 0),
      noblock_obuf_4_2_pipe_read_req => noblock_obuf_4_2_pipe_read_req(0 downto 0),
      noblock_obuf_4_2_pipe_read_ack => noblock_obuf_4_2_pipe_read_ack(0 downto 0),
      noblock_obuf_4_2_pipe_read_data => noblock_obuf_4_2_pipe_read_data(32 downto 0),
      noblock_obuf_2_2_pipe_read_req => noblock_obuf_2_2_pipe_read_req(0 downto 0),
      noblock_obuf_2_2_pipe_read_ack => noblock_obuf_2_2_pipe_read_ack(0 downto 0),
      noblock_obuf_2_2_pipe_read_data => noblock_obuf_2_2_pipe_read_data(32 downto 0),
      out_data_2_pipe_write_req => out_data_2_pipe_write_req(0 downto 0),
      out_data_2_pipe_write_ack => out_data_2_pipe_write_ack(0 downto 0),
      out_data_2_pipe_write_data => out_data_2_pipe_write_data(31 downto 0),
      updateCounter_call_reqs => updateCounter_call_reqs(3 downto 3),
      updateCounter_call_acks => updateCounter_call_acks(3 downto 3),
      updateCounter_call_data => updateCounter_call_data(67 downto 51),
      updateCounter_call_tag => updateCounter_call_tag(3 downto 3),
      updateCounter_return_reqs => updateCounter_return_reqs(3 downto 3),
      updateCounter_return_acks => updateCounter_return_acks(3 downto 3),
      updateCounter_return_data => updateCounter_return_data(3 downto 3),
      updateCounter_return_tag => updateCounter_return_tag(3 downto 3),
      tag_in => outputPort_2_Daemon_tag_in,
      tag_out => outputPort_2_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  outputPort_2_Daemon_tag_in <= (others => '0');
  outputPort_2_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => outputPort_2_Daemon_start_req, start_ack => outputPort_2_Daemon_start_ack,  fin_req => outputPort_2_Daemon_fin_req,  fin_ack => outputPort_2_Daemon_fin_ack);
  -- module outputPort_3_Daemon
  outputPort_3_Daemon_instance:outputPort_3_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => outputPort_3_Daemon_start_req,
      start_ack => outputPort_3_Daemon_start_ack,
      fin_req => outputPort_3_Daemon_fin_req,
      fin_ack => outputPort_3_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      noblock_obuf_1_3_pipe_read_req => noblock_obuf_1_3_pipe_read_req(0 downto 0),
      noblock_obuf_1_3_pipe_read_ack => noblock_obuf_1_3_pipe_read_ack(0 downto 0),
      noblock_obuf_1_3_pipe_read_data => noblock_obuf_1_3_pipe_read_data(32 downto 0),
      noblock_obuf_3_3_pipe_read_req => noblock_obuf_3_3_pipe_read_req(0 downto 0),
      noblock_obuf_3_3_pipe_read_ack => noblock_obuf_3_3_pipe_read_ack(0 downto 0),
      noblock_obuf_3_3_pipe_read_data => noblock_obuf_3_3_pipe_read_data(32 downto 0),
      noblock_obuf_4_3_pipe_read_req => noblock_obuf_4_3_pipe_read_req(0 downto 0),
      noblock_obuf_4_3_pipe_read_ack => noblock_obuf_4_3_pipe_read_ack(0 downto 0),
      noblock_obuf_4_3_pipe_read_data => noblock_obuf_4_3_pipe_read_data(32 downto 0),
      noblock_obuf_2_3_pipe_read_req => noblock_obuf_2_3_pipe_read_req(0 downto 0),
      noblock_obuf_2_3_pipe_read_ack => noblock_obuf_2_3_pipe_read_ack(0 downto 0),
      noblock_obuf_2_3_pipe_read_data => noblock_obuf_2_3_pipe_read_data(32 downto 0),
      out_data_3_pipe_write_req => out_data_3_pipe_write_req(0 downto 0),
      out_data_3_pipe_write_ack => out_data_3_pipe_write_ack(0 downto 0),
      out_data_3_pipe_write_data => out_data_3_pipe_write_data(31 downto 0),
      updateCounter_call_reqs => updateCounter_call_reqs(1 downto 1),
      updateCounter_call_acks => updateCounter_call_acks(1 downto 1),
      updateCounter_call_data => updateCounter_call_data(33 downto 17),
      updateCounter_call_tag => updateCounter_call_tag(1 downto 1),
      updateCounter_return_reqs => updateCounter_return_reqs(1 downto 1),
      updateCounter_return_acks => updateCounter_return_acks(1 downto 1),
      updateCounter_return_data => updateCounter_return_data(1 downto 1),
      updateCounter_return_tag => updateCounter_return_tag(1 downto 1),
      tag_in => outputPort_3_Daemon_tag_in,
      tag_out => outputPort_3_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  outputPort_3_Daemon_tag_in <= (others => '0');
  outputPort_3_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => outputPort_3_Daemon_start_req, start_ack => outputPort_3_Daemon_start_ack,  fin_req => outputPort_3_Daemon_fin_req,  fin_ack => outputPort_3_Daemon_fin_ack);
  -- module outputPort_4_Daemon
  outputPort_4_Daemon_instance:outputPort_4_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => outputPort_4_Daemon_start_req,
      start_ack => outputPort_4_Daemon_start_ack,
      fin_req => outputPort_4_Daemon_fin_req,
      fin_ack => outputPort_4_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      noblock_obuf_1_4_pipe_read_req => noblock_obuf_1_4_pipe_read_req(0 downto 0),
      noblock_obuf_1_4_pipe_read_ack => noblock_obuf_1_4_pipe_read_ack(0 downto 0),
      noblock_obuf_1_4_pipe_read_data => noblock_obuf_1_4_pipe_read_data(32 downto 0),
      noblock_obuf_3_4_pipe_read_req => noblock_obuf_3_4_pipe_read_req(0 downto 0),
      noblock_obuf_3_4_pipe_read_ack => noblock_obuf_3_4_pipe_read_ack(0 downto 0),
      noblock_obuf_3_4_pipe_read_data => noblock_obuf_3_4_pipe_read_data(32 downto 0),
      noblock_obuf_2_4_pipe_read_req => noblock_obuf_2_4_pipe_read_req(0 downto 0),
      noblock_obuf_2_4_pipe_read_ack => noblock_obuf_2_4_pipe_read_ack(0 downto 0),
      noblock_obuf_2_4_pipe_read_data => noblock_obuf_2_4_pipe_read_data(32 downto 0),
      noblock_obuf_4_4_pipe_read_req => noblock_obuf_4_4_pipe_read_req(0 downto 0),
      noblock_obuf_4_4_pipe_read_ack => noblock_obuf_4_4_pipe_read_ack(0 downto 0),
      noblock_obuf_4_4_pipe_read_data => noblock_obuf_4_4_pipe_read_data(32 downto 0),
      out_data_4_pipe_write_req => out_data_4_pipe_write_req(0 downto 0),
      out_data_4_pipe_write_ack => out_data_4_pipe_write_ack(0 downto 0),
      out_data_4_pipe_write_data => out_data_4_pipe_write_data(31 downto 0),
      updateCounter_call_reqs => updateCounter_call_reqs(0 downto 0),
      updateCounter_call_acks => updateCounter_call_acks(0 downto 0),
      updateCounter_call_data => updateCounter_call_data(16 downto 0),
      updateCounter_call_tag => updateCounter_call_tag(0 downto 0),
      updateCounter_return_reqs => updateCounter_return_reqs(0 downto 0),
      updateCounter_return_acks => updateCounter_return_acks(0 downto 0),
      updateCounter_return_data => updateCounter_return_data(0 downto 0),
      updateCounter_return_tag => updateCounter_return_tag(0 downto 0),
      tag_in => outputPort_4_Daemon_tag_in,
      tag_out => outputPort_4_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  outputPort_4_Daemon_tag_in <= (others => '0');
  outputPort_4_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => outputPort_4_Daemon_start_req, start_ack => outputPort_4_Daemon_start_ack,  fin_req => outputPort_4_Daemon_fin_req,  fin_ack => outputPort_4_Daemon_fin_ack);
  -- module updateCounter
  updateCounter_input_port <= updateCounter_in_args(16 downto 9);
  updateCounter_output_port <= updateCounter_in_args(8 downto 1);
  updateCounter_up <= updateCounter_in_args(0 downto 0);
  updateCounter_out_args <= updateCounter_continue ;
  -- call arbiter for module updateCounter
  updateCounter_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 8,
      call_data_width => 17,
      return_data_width => 1,
      callee_tag_length => 4,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => updateCounter_call_reqs,
      call_acks => updateCounter_call_acks,
      return_reqs => updateCounter_return_reqs,
      return_acks => updateCounter_return_acks,
      call_data  => updateCounter_call_data,
      call_tag  => updateCounter_call_tag,
      return_tag  => updateCounter_return_tag,
      call_mtag => updateCounter_tag_in,
      return_mtag => updateCounter_tag_out,
      return_data =>updateCounter_return_data,
      call_mreq => updateCounter_start_req,
      call_mack => updateCounter_start_ack,
      return_mreq => updateCounter_fin_req,
      return_mack => updateCounter_fin_ack,
      call_mdata => updateCounter_in_args,
      return_mdata => updateCounter_out_args,
      clk => clk, 
      reset => reset --
    ); --
  updateCounter_instance:updateCounter-- 
    generic map(tag_length => 5)
    port map(-- 
      input_port => updateCounter_input_port,
      output_port => updateCounter_output_port,
      up => updateCounter_up,
      continue => updateCounter_continue,
      start_req => updateCounter_start_req,
      start_ack => updateCounter_start_ack,
      fin_req => updateCounter_fin_req,
      fin_ack => updateCounter_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(3 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(19 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(1 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(2 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(3 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(1 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(19 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(2 downto 0),
      tag_in => updateCounter_tag_in,
      tag_out => updateCounter_tag_out-- 
    ); -- 
  in_data_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe in_data_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => in_data_1_pipe_read_req,
      read_ack => in_data_1_pipe_read_ack,
      read_data => in_data_1_pipe_read_data,
      write_req => in_data_1_pipe_write_req,
      write_ack => in_data_1_pipe_write_ack,
      write_data => in_data_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  in_data_2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe in_data_2",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => in_data_2_pipe_read_req,
      read_ack => in_data_2_pipe_read_ack,
      read_data => in_data_2_pipe_read_data,
      write_req => in_data_2_pipe_write_req,
      write_ack => in_data_2_pipe_write_ack,
      write_data => in_data_2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  in_data_3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe in_data_3",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => in_data_3_pipe_read_req,
      read_ack => in_data_3_pipe_read_ack,
      read_data => in_data_3_pipe_read_data,
      write_req => in_data_3_pipe_write_req,
      write_ack => in_data_3_pipe_write_ack,
      write_data => in_data_3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  in_data_4_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe in_data_4",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => in_data_4_pipe_read_req,
      read_ack => in_data_4_pipe_read_ack,
      read_data => in_data_4_pipe_read_data,
      write_req => in_data_4_pipe_write_req,
      write_ack => in_data_4_pipe_write_ack,
      write_data => in_data_4_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_1_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_1_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 128 --
    )
    port map( -- 
      read_req => noblock_obuf_1_1_pipe_read_req,
      read_ack => noblock_obuf_1_1_pipe_read_ack,
      read_data => noblock_obuf_1_1_pipe_read_data,
      write_req => noblock_obuf_1_1_pipe_write_req,
      write_ack => noblock_obuf_1_1_pipe_write_ack,
      write_data => noblock_obuf_1_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_1_2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_1_2",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 128 --
    )
    port map( -- 
      read_req => noblock_obuf_1_2_pipe_read_req,
      read_ack => noblock_obuf_1_2_pipe_read_ack,
      read_data => noblock_obuf_1_2_pipe_read_data,
      write_req => noblock_obuf_1_2_pipe_write_req,
      write_ack => noblock_obuf_1_2_pipe_write_ack,
      write_data => noblock_obuf_1_2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_1_3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_1_3",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 128 --
    )
    port map( -- 
      read_req => noblock_obuf_1_3_pipe_read_req,
      read_ack => noblock_obuf_1_3_pipe_read_ack,
      read_data => noblock_obuf_1_3_pipe_read_data,
      write_req => noblock_obuf_1_3_pipe_write_req,
      write_ack => noblock_obuf_1_3_pipe_write_ack,
      write_data => noblock_obuf_1_3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_1_4_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_1_4",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 128 --
    )
    port map( -- 
      read_req => noblock_obuf_1_4_pipe_read_req,
      read_ack => noblock_obuf_1_4_pipe_read_ack,
      read_data => noblock_obuf_1_4_pipe_read_data,
      write_req => noblock_obuf_1_4_pipe_write_req,
      write_ack => noblock_obuf_1_4_pipe_write_ack,
      write_data => noblock_obuf_1_4_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_2_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_2_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 128 --
    )
    port map( -- 
      read_req => noblock_obuf_2_1_pipe_read_req,
      read_ack => noblock_obuf_2_1_pipe_read_ack,
      read_data => noblock_obuf_2_1_pipe_read_data,
      write_req => noblock_obuf_2_1_pipe_write_req,
      write_ack => noblock_obuf_2_1_pipe_write_ack,
      write_data => noblock_obuf_2_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_2_2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_2_2",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 128 --
    )
    port map( -- 
      read_req => noblock_obuf_2_2_pipe_read_req,
      read_ack => noblock_obuf_2_2_pipe_read_ack,
      read_data => noblock_obuf_2_2_pipe_read_data,
      write_req => noblock_obuf_2_2_pipe_write_req,
      write_ack => noblock_obuf_2_2_pipe_write_ack,
      write_data => noblock_obuf_2_2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_2_3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_2_3",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 128 --
    )
    port map( -- 
      read_req => noblock_obuf_2_3_pipe_read_req,
      read_ack => noblock_obuf_2_3_pipe_read_ack,
      read_data => noblock_obuf_2_3_pipe_read_data,
      write_req => noblock_obuf_2_3_pipe_write_req,
      write_ack => noblock_obuf_2_3_pipe_write_ack,
      write_data => noblock_obuf_2_3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_2_4_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_2_4",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 128 --
    )
    port map( -- 
      read_req => noblock_obuf_2_4_pipe_read_req,
      read_ack => noblock_obuf_2_4_pipe_read_ack,
      read_data => noblock_obuf_2_4_pipe_read_data,
      write_req => noblock_obuf_2_4_pipe_write_req,
      write_ack => noblock_obuf_2_4_pipe_write_ack,
      write_data => noblock_obuf_2_4_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_3_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_3_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 128 --
    )
    port map( -- 
      read_req => noblock_obuf_3_1_pipe_read_req,
      read_ack => noblock_obuf_3_1_pipe_read_ack,
      read_data => noblock_obuf_3_1_pipe_read_data,
      write_req => noblock_obuf_3_1_pipe_write_req,
      write_ack => noblock_obuf_3_1_pipe_write_ack,
      write_data => noblock_obuf_3_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_3_2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_3_2",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 128 --
    )
    port map( -- 
      read_req => noblock_obuf_3_2_pipe_read_req,
      read_ack => noblock_obuf_3_2_pipe_read_ack,
      read_data => noblock_obuf_3_2_pipe_read_data,
      write_req => noblock_obuf_3_2_pipe_write_req,
      write_ack => noblock_obuf_3_2_pipe_write_ack,
      write_data => noblock_obuf_3_2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_3_3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_3_3",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 128 --
    )
    port map( -- 
      read_req => noblock_obuf_3_3_pipe_read_req,
      read_ack => noblock_obuf_3_3_pipe_read_ack,
      read_data => noblock_obuf_3_3_pipe_read_data,
      write_req => noblock_obuf_3_3_pipe_write_req,
      write_ack => noblock_obuf_3_3_pipe_write_ack,
      write_data => noblock_obuf_3_3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_3_4_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_3_4",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 128 --
    )
    port map( -- 
      read_req => noblock_obuf_3_4_pipe_read_req,
      read_ack => noblock_obuf_3_4_pipe_read_ack,
      read_data => noblock_obuf_3_4_pipe_read_data,
      write_req => noblock_obuf_3_4_pipe_write_req,
      write_ack => noblock_obuf_3_4_pipe_write_ack,
      write_data => noblock_obuf_3_4_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_4_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_4_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 128 --
    )
    port map( -- 
      read_req => noblock_obuf_4_1_pipe_read_req,
      read_ack => noblock_obuf_4_1_pipe_read_ack,
      read_data => noblock_obuf_4_1_pipe_read_data,
      write_req => noblock_obuf_4_1_pipe_write_req,
      write_ack => noblock_obuf_4_1_pipe_write_ack,
      write_data => noblock_obuf_4_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_4_2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_4_2",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 128 --
    )
    port map( -- 
      read_req => noblock_obuf_4_2_pipe_read_req,
      read_ack => noblock_obuf_4_2_pipe_read_ack,
      read_data => noblock_obuf_4_2_pipe_read_data,
      write_req => noblock_obuf_4_2_pipe_write_req,
      write_ack => noblock_obuf_4_2_pipe_write_ack,
      write_data => noblock_obuf_4_2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_4_3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_4_3",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 128 --
    )
    port map( -- 
      read_req => noblock_obuf_4_3_pipe_read_req,
      read_ack => noblock_obuf_4_3_pipe_read_ack,
      read_data => noblock_obuf_4_3_pipe_read_data,
      write_req => noblock_obuf_4_3_pipe_write_req,
      write_ack => noblock_obuf_4_3_pipe_write_ack,
      write_data => noblock_obuf_4_3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_4_4_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_4_4",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 128 --
    )
    port map( -- 
      read_req => noblock_obuf_4_4_pipe_read_req,
      read_ack => noblock_obuf_4_4_pipe_read_ack,
      read_data => noblock_obuf_4_4_pipe_read_data,
      write_req => noblock_obuf_4_4_pipe_write_req,
      write_ack => noblock_obuf_4_4_pipe_write_ack,
      write_data => noblock_obuf_4_4_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_data_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe out_data_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => out_data_1_pipe_read_req,
      read_ack => out_data_1_pipe_read_ack,
      read_data => out_data_1_pipe_read_data,
      write_req => out_data_1_pipe_write_req,
      write_ack => out_data_1_pipe_write_ack,
      write_data => out_data_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_data_2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe out_data_2",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => out_data_2_pipe_read_req,
      read_ack => out_data_2_pipe_read_ack,
      read_data => out_data_2_pipe_read_data,
      write_req => out_data_2_pipe_write_req,
      write_ack => out_data_2_pipe_write_ack,
      write_data => out_data_2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_data_3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe out_data_3",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => out_data_3_pipe_read_req,
      read_ack => out_data_3_pipe_read_ack,
      read_data => out_data_3_pipe_read_data,
      write_req => out_data_3_pipe_write_req,
      write_ack => out_data_3_pipe_write_ack,
      write_data => out_data_3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_data_4_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe out_data_4",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => out_data_4_pipe_read_req,
      read_ack => out_data_4_pipe_read_ack,
      read_data => out_data_4_pipe_read_data,
      write_req => out_data_4_pipe_write_req,
      write_ack => out_data_4_pipe_write_ack,
      write_data => out_data_4_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 2,
      addr_width => 4,
      data_width => 2,
      tag_width => 3,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 4,
      base_bank_data_width => 2
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
